module MG_FA(
  input a,
  input b,
  input cin,
  output sum,
  output cout
);

  assign sum = (a ^ b) ^ cin;
  assign cout = (a & b) | (b & cin) | (a & cin);
endmodule
module MG_HA(
  input a,
  input b,
  output sum,
  output cout
);

  assign sum = a ^ b;
  assign cout = a & b;
endmodule
module mult16s_normal_brentkung(
  input [15:0] multiplicand,
  input [15:0] multiplier,
  output [31:0] product
);

  wire pp_0_0;
  wire pp_0_1;
  wire pp_0_10;
  wire pp_0_11;
  wire pp_0_12;
  wire pp_0_13;
  wire pp_0_14;
  wire pp_0_15;
  wire pp_0_16;
  wire pp_0_2;
  wire pp_0_3;
  wire pp_0_4;
  wire pp_0_5;
  wire pp_0_6;
  wire pp_0_7;
  wire pp_0_8;
  wire pp_0_9;
  wire pp_10_10;
  wire pp_10_11;
  wire pp_10_12;
  wire pp_10_13;
  wire pp_10_14;
  wire pp_10_15;
  wire pp_10_16;
  wire pp_10_17;
  wire pp_10_18;
  wire pp_10_19;
  wire pp_10_20;
  wire pp_10_21;
  wire pp_10_22;
  wire pp_10_23;
  wire pp_10_24;
  wire pp_10_25;
  wire pp_11_11;
  wire pp_11_12;
  wire pp_11_13;
  wire pp_11_14;
  wire pp_11_15;
  wire pp_11_16;
  wire pp_11_17;
  wire pp_11_18;
  wire pp_11_19;
  wire pp_11_20;
  wire pp_11_21;
  wire pp_11_22;
  wire pp_11_23;
  wire pp_11_24;
  wire pp_11_25;
  wire pp_11_26;
  wire pp_12_12;
  wire pp_12_13;
  wire pp_12_14;
  wire pp_12_15;
  wire pp_12_16;
  wire pp_12_17;
  wire pp_12_18;
  wire pp_12_19;
  wire pp_12_20;
  wire pp_12_21;
  wire pp_12_22;
  wire pp_12_23;
  wire pp_12_24;
  wire pp_12_25;
  wire pp_12_26;
  wire pp_12_27;
  wire pp_13_13;
  wire pp_13_14;
  wire pp_13_15;
  wire pp_13_16;
  wire pp_13_17;
  wire pp_13_18;
  wire pp_13_19;
  wire pp_13_20;
  wire pp_13_21;
  wire pp_13_22;
  wire pp_13_23;
  wire pp_13_24;
  wire pp_13_25;
  wire pp_13_26;
  wire pp_13_27;
  wire pp_13_28;
  wire pp_14_14;
  wire pp_14_15;
  wire pp_14_16;
  wire pp_14_17;
  wire pp_14_18;
  wire pp_14_19;
  wire pp_14_20;
  wire pp_14_21;
  wire pp_14_22;
  wire pp_14_23;
  wire pp_14_24;
  wire pp_14_25;
  wire pp_14_26;
  wire pp_14_27;
  wire pp_14_28;
  wire pp_14_29;
  wire pp_15_15;
  wire pp_15_16;
  wire pp_15_17;
  wire pp_15_18;
  wire pp_15_19;
  wire pp_15_20;
  wire pp_15_21;
  wire pp_15_22;
  wire pp_15_23;
  wire pp_15_24;
  wire pp_15_25;
  wire pp_15_26;
  wire pp_15_27;
  wire pp_15_28;
  wire pp_15_29;
  wire pp_15_30;
  wire pp_15_31;
  wire pp_1_1;
  wire pp_1_10;
  wire pp_1_11;
  wire pp_1_12;
  wire pp_1_13;
  wire pp_1_14;
  wire pp_1_15;
  wire pp_1_16;
  wire pp_1_2;
  wire pp_1_3;
  wire pp_1_4;
  wire pp_1_5;
  wire pp_1_6;
  wire pp_1_7;
  wire pp_1_8;
  wire pp_1_9;
  wire pp_2_10;
  wire pp_2_11;
  wire pp_2_12;
  wire pp_2_13;
  wire pp_2_14;
  wire pp_2_15;
  wire pp_2_16;
  wire pp_2_17;
  wire pp_2_2;
  wire pp_2_3;
  wire pp_2_4;
  wire pp_2_5;
  wire pp_2_6;
  wire pp_2_7;
  wire pp_2_8;
  wire pp_2_9;
  wire pp_3_10;
  wire pp_3_11;
  wire pp_3_12;
  wire pp_3_13;
  wire pp_3_14;
  wire pp_3_15;
  wire pp_3_16;
  wire pp_3_17;
  wire pp_3_18;
  wire pp_3_3;
  wire pp_3_4;
  wire pp_3_5;
  wire pp_3_6;
  wire pp_3_7;
  wire pp_3_8;
  wire pp_3_9;
  wire pp_4_10;
  wire pp_4_11;
  wire pp_4_12;
  wire pp_4_13;
  wire pp_4_14;
  wire pp_4_15;
  wire pp_4_16;
  wire pp_4_17;
  wire pp_4_18;
  wire pp_4_19;
  wire pp_4_4;
  wire pp_4_5;
  wire pp_4_6;
  wire pp_4_7;
  wire pp_4_8;
  wire pp_4_9;
  wire pp_5_10;
  wire pp_5_11;
  wire pp_5_12;
  wire pp_5_13;
  wire pp_5_14;
  wire pp_5_15;
  wire pp_5_16;
  wire pp_5_17;
  wire pp_5_18;
  wire pp_5_19;
  wire pp_5_20;
  wire pp_5_5;
  wire pp_5_6;
  wire pp_5_7;
  wire pp_5_8;
  wire pp_5_9;
  wire pp_6_10;
  wire pp_6_11;
  wire pp_6_12;
  wire pp_6_13;
  wire pp_6_14;
  wire pp_6_15;
  wire pp_6_16;
  wire pp_6_17;
  wire pp_6_18;
  wire pp_6_19;
  wire pp_6_20;
  wire pp_6_21;
  wire pp_6_6;
  wire pp_6_7;
  wire pp_6_8;
  wire pp_6_9;
  wire pp_7_10;
  wire pp_7_11;
  wire pp_7_12;
  wire pp_7_13;
  wire pp_7_14;
  wire pp_7_15;
  wire pp_7_16;
  wire pp_7_17;
  wire pp_7_18;
  wire pp_7_19;
  wire pp_7_20;
  wire pp_7_21;
  wire pp_7_22;
  wire pp_7_7;
  wire pp_7_8;
  wire pp_7_9;
  wire pp_8_10;
  wire pp_8_11;
  wire pp_8_12;
  wire pp_8_13;
  wire pp_8_14;
  wire pp_8_15;
  wire pp_8_16;
  wire pp_8_17;
  wire pp_8_18;
  wire pp_8_19;
  wire pp_8_20;
  wire pp_8_21;
  wire pp_8_22;
  wire pp_8_23;
  wire pp_8_8;
  wire pp_8_9;
  wire pp_9_10;
  wire pp_9_11;
  wire pp_9_12;
  wire pp_9_13;
  wire pp_9_14;
  wire pp_9_15;
  wire pp_9_16;
  wire pp_9_17;
  wire pp_9_18;
  wire pp_9_19;
  wire pp_9_20;
  wire pp_9_21;
  wire pp_9_22;
  wire pp_9_23;
  wire pp_9_24;
  wire pp_9_9;
  assign pp_0_0 = multiplicand[0] & multiplier[0];
  assign pp_0_1 = multiplicand[1] & multiplier[0];
  assign pp_0_10 = multiplicand[10] & multiplier[0];
  assign pp_0_11 = multiplicand[11] & multiplier[0];
  assign pp_0_12 = multiplicand[12] & multiplier[0];
  assign pp_0_13 = multiplicand[13] & multiplier[0];
  assign pp_0_14 = multiplicand[14] & multiplier[0];
  assign pp_0_15 = ~(multiplicand[15] & multiplier[0]);
  assign pp_0_16 = multiplier[15];
  assign pp_0_2 = multiplicand[2] & multiplier[0];
  assign pp_0_3 = multiplicand[3] & multiplier[0];
  assign pp_0_4 = multiplicand[4] & multiplier[0];
  assign pp_0_5 = multiplicand[5] & multiplier[0];
  assign pp_0_6 = multiplicand[6] & multiplier[0];
  assign pp_0_7 = multiplicand[7] & multiplier[0];
  assign pp_0_8 = multiplicand[8] & multiplier[0];
  assign pp_0_9 = multiplicand[9] & multiplier[0];
  assign pp_10_10 = multiplicand[0] & multiplier[10];
  assign pp_10_11 = multiplicand[1] & multiplier[10];
  assign pp_10_12 = multiplicand[2] & multiplier[10];
  assign pp_10_13 = multiplicand[3] & multiplier[10];
  assign pp_10_14 = multiplicand[4] & multiplier[10];
  assign pp_10_15 = multiplicand[5] & multiplier[10];
  assign pp_10_16 = multiplicand[6] & multiplier[10];
  assign pp_10_17 = multiplicand[7] & multiplier[10];
  assign pp_10_18 = multiplicand[8] & multiplier[10];
  assign pp_10_19 = multiplicand[9] & multiplier[10];
  assign pp_10_20 = multiplicand[10] & multiplier[10];
  assign pp_10_21 = multiplicand[11] & multiplier[10];
  assign pp_10_22 = multiplicand[12] & multiplier[10];
  assign pp_10_23 = multiplicand[13] & multiplier[10];
  assign pp_10_24 = multiplicand[14] & multiplier[10];
  assign pp_10_25 = ~(multiplicand[15] & multiplier[10]);
  assign pp_11_11 = multiplicand[0] & multiplier[11];
  assign pp_11_12 = multiplicand[1] & multiplier[11];
  assign pp_11_13 = multiplicand[2] & multiplier[11];
  assign pp_11_14 = multiplicand[3] & multiplier[11];
  assign pp_11_15 = multiplicand[4] & multiplier[11];
  assign pp_11_16 = multiplicand[5] & multiplier[11];
  assign pp_11_17 = multiplicand[6] & multiplier[11];
  assign pp_11_18 = multiplicand[7] & multiplier[11];
  assign pp_11_19 = multiplicand[8] & multiplier[11];
  assign pp_11_20 = multiplicand[9] & multiplier[11];
  assign pp_11_21 = multiplicand[10] & multiplier[11];
  assign pp_11_22 = multiplicand[11] & multiplier[11];
  assign pp_11_23 = multiplicand[12] & multiplier[11];
  assign pp_11_24 = multiplicand[13] & multiplier[11];
  assign pp_11_25 = multiplicand[14] & multiplier[11];
  assign pp_11_26 = ~(multiplicand[15] & multiplier[11]);
  assign pp_12_12 = multiplicand[0] & multiplier[12];
  assign pp_12_13 = multiplicand[1] & multiplier[12];
  assign pp_12_14 = multiplicand[2] & multiplier[12];
  assign pp_12_15 = multiplicand[3] & multiplier[12];
  assign pp_12_16 = multiplicand[4] & multiplier[12];
  assign pp_12_17 = multiplicand[5] & multiplier[12];
  assign pp_12_18 = multiplicand[6] & multiplier[12];
  assign pp_12_19 = multiplicand[7] & multiplier[12];
  assign pp_12_20 = multiplicand[8] & multiplier[12];
  assign pp_12_21 = multiplicand[9] & multiplier[12];
  assign pp_12_22 = multiplicand[10] & multiplier[12];
  assign pp_12_23 = multiplicand[11] & multiplier[12];
  assign pp_12_24 = multiplicand[12] & multiplier[12];
  assign pp_12_25 = multiplicand[13] & multiplier[12];
  assign pp_12_26 = multiplicand[14] & multiplier[12];
  assign pp_12_27 = ~(multiplicand[15] & multiplier[12]);
  assign pp_13_13 = multiplicand[0] & multiplier[13];
  assign pp_13_14 = multiplicand[1] & multiplier[13];
  assign pp_13_15 = multiplicand[2] & multiplier[13];
  assign pp_13_16 = multiplicand[3] & multiplier[13];
  assign pp_13_17 = multiplicand[4] & multiplier[13];
  assign pp_13_18 = multiplicand[5] & multiplier[13];
  assign pp_13_19 = multiplicand[6] & multiplier[13];
  assign pp_13_20 = multiplicand[7] & multiplier[13];
  assign pp_13_21 = multiplicand[8] & multiplier[13];
  assign pp_13_22 = multiplicand[9] & multiplier[13];
  assign pp_13_23 = multiplicand[10] & multiplier[13];
  assign pp_13_24 = multiplicand[11] & multiplier[13];
  assign pp_13_25 = multiplicand[12] & multiplier[13];
  assign pp_13_26 = multiplicand[13] & multiplier[13];
  assign pp_13_27 = multiplicand[14] & multiplier[13];
  assign pp_13_28 = ~(multiplicand[15] & multiplier[13]);
  assign pp_14_14 = multiplicand[0] & multiplier[14];
  assign pp_14_15 = multiplicand[1] & multiplier[14];
  assign pp_14_16 = multiplicand[2] & multiplier[14];
  assign pp_14_17 = multiplicand[3] & multiplier[14];
  assign pp_14_18 = multiplicand[4] & multiplier[14];
  assign pp_14_19 = multiplicand[5] & multiplier[14];
  assign pp_14_20 = multiplicand[6] & multiplier[14];
  assign pp_14_21 = multiplicand[7] & multiplier[14];
  assign pp_14_22 = multiplicand[8] & multiplier[14];
  assign pp_14_23 = multiplicand[9] & multiplier[14];
  assign pp_14_24 = multiplicand[10] & multiplier[14];
  assign pp_14_25 = multiplicand[11] & multiplier[14];
  assign pp_14_26 = multiplicand[12] & multiplier[14];
  assign pp_14_27 = multiplicand[13] & multiplier[14];
  assign pp_14_28 = multiplicand[14] & multiplier[14];
  assign pp_14_29 = ~(multiplicand[15] & multiplier[14]);
  assign pp_15_15 = ~(multiplicand[0] & multiplier[15]);
  assign pp_15_16 = ~multiplicand[1] & multiplier[15];
  assign pp_15_17 = ~multiplicand[2] & multiplier[15];
  assign pp_15_18 = ~multiplicand[3] & multiplier[15];
  assign pp_15_19 = ~multiplicand[4] & multiplier[15];
  assign pp_15_20 = ~multiplicand[5] & multiplier[15];
  assign pp_15_21 = ~multiplicand[6] & multiplier[15];
  assign pp_15_22 = ~multiplicand[7] & multiplier[15];
  assign pp_15_23 = ~multiplicand[8] & multiplier[15];
  assign pp_15_24 = ~multiplicand[9] & multiplier[15];
  assign pp_15_25 = ~multiplicand[10] & multiplier[15];
  assign pp_15_26 = ~multiplicand[11] & multiplier[15];
  assign pp_15_27 = ~multiplicand[12] & multiplier[15];
  assign pp_15_28 = ~multiplicand[13] & multiplier[15];
  assign pp_15_29 = ~multiplicand[14] & multiplier[15];
  assign pp_15_30 = ~(~multiplicand[15] & multiplier[15]);
  assign pp_15_31 = 1'b1;
  assign pp_1_1 = multiplicand[0] & multiplier[1];
  assign pp_1_10 = multiplicand[9] & multiplier[1];
  assign pp_1_11 = multiplicand[10] & multiplier[1];
  assign pp_1_12 = multiplicand[11] & multiplier[1];
  assign pp_1_13 = multiplicand[12] & multiplier[1];
  assign pp_1_14 = multiplicand[13] & multiplier[1];
  assign pp_1_15 = multiplicand[14] & multiplier[1];
  assign pp_1_16 = ~(multiplicand[15] & multiplier[1]);
  assign pp_1_2 = multiplicand[1] & multiplier[1];
  assign pp_1_3 = multiplicand[2] & multiplier[1];
  assign pp_1_4 = multiplicand[3] & multiplier[1];
  assign pp_1_5 = multiplicand[4] & multiplier[1];
  assign pp_1_6 = multiplicand[5] & multiplier[1];
  assign pp_1_7 = multiplicand[6] & multiplier[1];
  assign pp_1_8 = multiplicand[7] & multiplier[1];
  assign pp_1_9 = multiplicand[8] & multiplier[1];
  assign pp_2_10 = multiplicand[8] & multiplier[2];
  assign pp_2_11 = multiplicand[9] & multiplier[2];
  assign pp_2_12 = multiplicand[10] & multiplier[2];
  assign pp_2_13 = multiplicand[11] & multiplier[2];
  assign pp_2_14 = multiplicand[12] & multiplier[2];
  assign pp_2_15 = multiplicand[13] & multiplier[2];
  assign pp_2_16 = multiplicand[14] & multiplier[2];
  assign pp_2_17 = ~(multiplicand[15] & multiplier[2]);
  assign pp_2_2 = multiplicand[0] & multiplier[2];
  assign pp_2_3 = multiplicand[1] & multiplier[2];
  assign pp_2_4 = multiplicand[2] & multiplier[2];
  assign pp_2_5 = multiplicand[3] & multiplier[2];
  assign pp_2_6 = multiplicand[4] & multiplier[2];
  assign pp_2_7 = multiplicand[5] & multiplier[2];
  assign pp_2_8 = multiplicand[6] & multiplier[2];
  assign pp_2_9 = multiplicand[7] & multiplier[2];
  assign pp_3_10 = multiplicand[7] & multiplier[3];
  assign pp_3_11 = multiplicand[8] & multiplier[3];
  assign pp_3_12 = multiplicand[9] & multiplier[3];
  assign pp_3_13 = multiplicand[10] & multiplier[3];
  assign pp_3_14 = multiplicand[11] & multiplier[3];
  assign pp_3_15 = multiplicand[12] & multiplier[3];
  assign pp_3_16 = multiplicand[13] & multiplier[3];
  assign pp_3_17 = multiplicand[14] & multiplier[3];
  assign pp_3_18 = ~(multiplicand[15] & multiplier[3]);
  assign pp_3_3 = multiplicand[0] & multiplier[3];
  assign pp_3_4 = multiplicand[1] & multiplier[3];
  assign pp_3_5 = multiplicand[2] & multiplier[3];
  assign pp_3_6 = multiplicand[3] & multiplier[3];
  assign pp_3_7 = multiplicand[4] & multiplier[3];
  assign pp_3_8 = multiplicand[5] & multiplier[3];
  assign pp_3_9 = multiplicand[6] & multiplier[3];
  assign pp_4_10 = multiplicand[6] & multiplier[4];
  assign pp_4_11 = multiplicand[7] & multiplier[4];
  assign pp_4_12 = multiplicand[8] & multiplier[4];
  assign pp_4_13 = multiplicand[9] & multiplier[4];
  assign pp_4_14 = multiplicand[10] & multiplier[4];
  assign pp_4_15 = multiplicand[11] & multiplier[4];
  assign pp_4_16 = multiplicand[12] & multiplier[4];
  assign pp_4_17 = multiplicand[13] & multiplier[4];
  assign pp_4_18 = multiplicand[14] & multiplier[4];
  assign pp_4_19 = ~(multiplicand[15] & multiplier[4]);
  assign pp_4_4 = multiplicand[0] & multiplier[4];
  assign pp_4_5 = multiplicand[1] & multiplier[4];
  assign pp_4_6 = multiplicand[2] & multiplier[4];
  assign pp_4_7 = multiplicand[3] & multiplier[4];
  assign pp_4_8 = multiplicand[4] & multiplier[4];
  assign pp_4_9 = multiplicand[5] & multiplier[4];
  assign pp_5_10 = multiplicand[5] & multiplier[5];
  assign pp_5_11 = multiplicand[6] & multiplier[5];
  assign pp_5_12 = multiplicand[7] & multiplier[5];
  assign pp_5_13 = multiplicand[8] & multiplier[5];
  assign pp_5_14 = multiplicand[9] & multiplier[5];
  assign pp_5_15 = multiplicand[10] & multiplier[5];
  assign pp_5_16 = multiplicand[11] & multiplier[5];
  assign pp_5_17 = multiplicand[12] & multiplier[5];
  assign pp_5_18 = multiplicand[13] & multiplier[5];
  assign pp_5_19 = multiplicand[14] & multiplier[5];
  assign pp_5_20 = ~(multiplicand[15] & multiplier[5]);
  assign pp_5_5 = multiplicand[0] & multiplier[5];
  assign pp_5_6 = multiplicand[1] & multiplier[5];
  assign pp_5_7 = multiplicand[2] & multiplier[5];
  assign pp_5_8 = multiplicand[3] & multiplier[5];
  assign pp_5_9 = multiplicand[4] & multiplier[5];
  assign pp_6_10 = multiplicand[4] & multiplier[6];
  assign pp_6_11 = multiplicand[5] & multiplier[6];
  assign pp_6_12 = multiplicand[6] & multiplier[6];
  assign pp_6_13 = multiplicand[7] & multiplier[6];
  assign pp_6_14 = multiplicand[8] & multiplier[6];
  assign pp_6_15 = multiplicand[9] & multiplier[6];
  assign pp_6_16 = multiplicand[10] & multiplier[6];
  assign pp_6_17 = multiplicand[11] & multiplier[6];
  assign pp_6_18 = multiplicand[12] & multiplier[6];
  assign pp_6_19 = multiplicand[13] & multiplier[6];
  assign pp_6_20 = multiplicand[14] & multiplier[6];
  assign pp_6_21 = ~(multiplicand[15] & multiplier[6]);
  assign pp_6_6 = multiplicand[0] & multiplier[6];
  assign pp_6_7 = multiplicand[1] & multiplier[6];
  assign pp_6_8 = multiplicand[2] & multiplier[6];
  assign pp_6_9 = multiplicand[3] & multiplier[6];
  assign pp_7_10 = multiplicand[3] & multiplier[7];
  assign pp_7_11 = multiplicand[4] & multiplier[7];
  assign pp_7_12 = multiplicand[5] & multiplier[7];
  assign pp_7_13 = multiplicand[6] & multiplier[7];
  assign pp_7_14 = multiplicand[7] & multiplier[7];
  assign pp_7_15 = multiplicand[8] & multiplier[7];
  assign pp_7_16 = multiplicand[9] & multiplier[7];
  assign pp_7_17 = multiplicand[10] & multiplier[7];
  assign pp_7_18 = multiplicand[11] & multiplier[7];
  assign pp_7_19 = multiplicand[12] & multiplier[7];
  assign pp_7_20 = multiplicand[13] & multiplier[7];
  assign pp_7_21 = multiplicand[14] & multiplier[7];
  assign pp_7_22 = ~(multiplicand[15] & multiplier[7]);
  assign pp_7_7 = multiplicand[0] & multiplier[7];
  assign pp_7_8 = multiplicand[1] & multiplier[7];
  assign pp_7_9 = multiplicand[2] & multiplier[7];
  assign pp_8_10 = multiplicand[2] & multiplier[8];
  assign pp_8_11 = multiplicand[3] & multiplier[8];
  assign pp_8_12 = multiplicand[4] & multiplier[8];
  assign pp_8_13 = multiplicand[5] & multiplier[8];
  assign pp_8_14 = multiplicand[6] & multiplier[8];
  assign pp_8_15 = multiplicand[7] & multiplier[8];
  assign pp_8_16 = multiplicand[8] & multiplier[8];
  assign pp_8_17 = multiplicand[9] & multiplier[8];
  assign pp_8_18 = multiplicand[10] & multiplier[8];
  assign pp_8_19 = multiplicand[11] & multiplier[8];
  assign pp_8_20 = multiplicand[12] & multiplier[8];
  assign pp_8_21 = multiplicand[13] & multiplier[8];
  assign pp_8_22 = multiplicand[14] & multiplier[8];
  assign pp_8_23 = ~(multiplicand[15] & multiplier[8]);
  assign pp_8_8 = multiplicand[0] & multiplier[8];
  assign pp_8_9 = multiplicand[1] & multiplier[8];
  assign pp_9_10 = multiplicand[1] & multiplier[9];
  assign pp_9_11 = multiplicand[2] & multiplier[9];
  assign pp_9_12 = multiplicand[3] & multiplier[9];
  assign pp_9_13 = multiplicand[4] & multiplier[9];
  assign pp_9_14 = multiplicand[5] & multiplier[9];
  assign pp_9_15 = multiplicand[6] & multiplier[9];
  assign pp_9_16 = multiplicand[7] & multiplier[9];
  assign pp_9_17 = multiplicand[8] & multiplier[9];
  assign pp_9_18 = multiplicand[9] & multiplier[9];
  assign pp_9_19 = multiplicand[10] & multiplier[9];
  assign pp_9_20 = multiplicand[11] & multiplier[9];
  assign pp_9_21 = multiplicand[12] & multiplier[9];
  assign pp_9_22 = multiplicand[13] & multiplier[9];
  assign pp_9_23 = multiplicand[14] & multiplier[9];
  assign pp_9_24 = ~(multiplicand[15] & multiplier[9]);
  assign pp_9_9 = multiplicand[0] & multiplier[9];
  wire pp_0_0_0;
  wire pp_0_1_0;
  wire pp_0_1_1;
  wire pp_0_2_0;
  wire pp_0_2_1;
  wire pp_0_2_2;
  wire pp_0_3_0;
  wire pp_0_3_1;
  wire pp_0_3_2;
  wire pp_0_3_3;
  wire pp_0_4_0;
  wire pp_0_4_1;
  wire pp_0_4_2;
  wire pp_0_4_3;
  wire pp_0_4_4;
  wire pp_0_5_0;
  wire pp_0_5_1;
  wire pp_0_5_2;
  wire pp_0_5_3;
  wire pp_0_5_4;
  wire pp_0_5_5;
  wire pp_0_6_0;
  wire pp_0_6_1;
  wire pp_0_6_2;
  wire pp_0_6_3;
  wire pp_0_6_4;
  wire pp_0_6_5;
  wire pp_0_6_6;
  wire pp_0_7_0;
  wire pp_0_7_1;
  wire pp_0_7_2;
  wire pp_0_7_3;
  wire pp_0_7_4;
  wire pp_0_7_5;
  wire pp_0_7_6;
  wire pp_0_7_7;
  wire pp_0_8_0;
  wire pp_0_8_1;
  wire pp_0_8_2;
  wire pp_0_8_3;
  wire pp_0_8_4;
  wire pp_0_8_5;
  wire pp_0_8_6;
  wire pp_0_8_7;
  wire pp_0_8_8;
  wire pp_0_9_0;
  wire pp_0_9_1;
  wire pp_0_9_2;
  wire pp_0_9_3;
  wire pp_0_9_4;
  wire pp_0_9_5;
  wire pp_0_9_6;
  wire pp_0_9_7;
  wire pp_0_9_8;
  wire pp_0_9_9;
  wire pp_0_10_0;
  wire pp_0_10_1;
  wire pp_0_10_2;
  wire pp_0_10_3;
  wire pp_0_10_4;
  wire pp_0_10_5;
  wire pp_0_10_6;
  wire pp_0_10_7;
  wire pp_0_10_8;
  wire pp_0_10_9;
  wire pp_0_10_10;
  wire pp_0_11_0;
  wire pp_0_11_1;
  wire pp_0_11_2;
  wire pp_0_11_3;
  wire pp_0_11_4;
  wire pp_0_11_5;
  wire pp_0_11_6;
  wire pp_0_11_7;
  wire pp_0_11_8;
  wire pp_0_11_9;
  wire pp_0_11_10;
  wire pp_0_11_11;
  wire pp_0_12_0;
  wire pp_0_12_1;
  wire pp_0_12_2;
  wire pp_0_12_3;
  wire pp_0_12_4;
  wire pp_0_12_5;
  wire pp_0_12_6;
  wire pp_0_12_7;
  wire pp_0_12_8;
  wire pp_0_12_9;
  wire pp_0_12_10;
  wire pp_0_12_11;
  wire pp_0_12_12;
  wire pp_0_13_0;
  wire pp_0_13_1;
  wire pp_0_13_2;
  wire pp_0_13_3;
  wire pp_0_13_4;
  wire pp_0_13_5;
  wire pp_0_13_6;
  wire pp_0_13_7;
  wire pp_0_13_8;
  wire pp_0_13_9;
  wire pp_0_13_10;
  wire pp_0_13_11;
  wire pp_0_13_12;
  wire pp_0_13_13;
  wire pp_0_14_0;
  wire pp_0_14_1;
  wire pp_0_14_2;
  wire pp_0_14_3;
  wire pp_0_14_4;
  wire pp_0_14_5;
  wire pp_0_14_6;
  wire pp_0_14_7;
  wire pp_0_14_8;
  wire pp_0_14_9;
  wire pp_0_14_10;
  wire pp_0_14_11;
  wire pp_0_14_12;
  wire pp_0_14_13;
  wire pp_0_14_14;
  wire pp_0_15_0;
  wire pp_0_15_1;
  wire pp_0_15_2;
  wire pp_0_15_3;
  wire pp_0_15_4;
  wire pp_0_15_5;
  wire pp_0_15_6;
  wire pp_0_15_7;
  wire pp_0_15_8;
  wire pp_0_15_9;
  wire pp_0_15_10;
  wire pp_0_15_11;
  wire pp_0_15_12;
  wire pp_0_15_13;
  wire pp_0_15_14;
  wire pp_0_15_15;
  wire pp_0_16_0;
  wire pp_0_16_1;
  wire pp_0_16_2;
  wire pp_0_16_3;
  wire pp_0_16_4;
  wire pp_0_16_5;
  wire pp_0_16_6;
  wire pp_0_16_7;
  wire pp_0_16_8;
  wire pp_0_16_9;
  wire pp_0_16_10;
  wire pp_0_16_11;
  wire pp_0_16_12;
  wire pp_0_16_13;
  wire pp_0_16_14;
  wire pp_0_16_15;
  wire pp_0_17_0;
  wire pp_0_17_1;
  wire pp_0_17_2;
  wire pp_0_17_3;
  wire pp_0_17_4;
  wire pp_0_17_5;
  wire pp_0_17_6;
  wire pp_0_17_7;
  wire pp_0_17_8;
  wire pp_0_17_9;
  wire pp_0_17_10;
  wire pp_0_17_11;
  wire pp_0_17_12;
  wire pp_0_17_13;
  wire pp_0_18_0;
  wire pp_0_18_1;
  wire pp_0_18_2;
  wire pp_0_18_3;
  wire pp_0_18_4;
  wire pp_0_18_5;
  wire pp_0_18_6;
  wire pp_0_18_7;
  wire pp_0_18_8;
  wire pp_0_18_9;
  wire pp_0_18_10;
  wire pp_0_18_11;
  wire pp_0_18_12;
  wire pp_0_19_0;
  wire pp_0_19_1;
  wire pp_0_19_2;
  wire pp_0_19_3;
  wire pp_0_19_4;
  wire pp_0_19_5;
  wire pp_0_19_6;
  wire pp_0_19_7;
  wire pp_0_19_8;
  wire pp_0_19_9;
  wire pp_0_19_10;
  wire pp_0_19_11;
  wire pp_0_20_0;
  wire pp_0_20_1;
  wire pp_0_20_2;
  wire pp_0_20_3;
  wire pp_0_20_4;
  wire pp_0_20_5;
  wire pp_0_20_6;
  wire pp_0_20_7;
  wire pp_0_20_8;
  wire pp_0_20_9;
  wire pp_0_20_10;
  wire pp_0_21_0;
  wire pp_0_21_1;
  wire pp_0_21_2;
  wire pp_0_21_3;
  wire pp_0_21_4;
  wire pp_0_21_5;
  wire pp_0_21_6;
  wire pp_0_21_7;
  wire pp_0_21_8;
  wire pp_0_21_9;
  wire pp_0_22_0;
  wire pp_0_22_1;
  wire pp_0_22_2;
  wire pp_0_22_3;
  wire pp_0_22_4;
  wire pp_0_22_5;
  wire pp_0_22_6;
  wire pp_0_22_7;
  wire pp_0_22_8;
  wire pp_0_23_0;
  wire pp_0_23_1;
  wire pp_0_23_2;
  wire pp_0_23_3;
  wire pp_0_23_4;
  wire pp_0_23_5;
  wire pp_0_23_6;
  wire pp_0_23_7;
  wire pp_0_24_0;
  wire pp_0_24_1;
  wire pp_0_24_2;
  wire pp_0_24_3;
  wire pp_0_24_4;
  wire pp_0_24_5;
  wire pp_0_24_6;
  wire pp_0_25_0;
  wire pp_0_25_1;
  wire pp_0_25_2;
  wire pp_0_25_3;
  wire pp_0_25_4;
  wire pp_0_25_5;
  wire pp_0_26_0;
  wire pp_0_26_1;
  wire pp_0_26_2;
  wire pp_0_26_3;
  wire pp_0_26_4;
  wire pp_0_27_0;
  wire pp_0_27_1;
  wire pp_0_27_2;
  wire pp_0_27_3;
  wire pp_0_28_0;
  wire pp_0_28_1;
  wire pp_0_28_2;
  wire pp_0_29_0;
  wire pp_0_29_1;
  wire pp_0_30_0;
  wire pp_0_31_0;
  wire pp_1_0_0;
  wire pp_1_1_0;
  wire pp_1_1_1;
  wire pp_1_2_0;
  wire pp_1_2_1;
  wire pp_1_2_2;
  wire pp_1_3_0;
  wire pp_1_3_1;
  wire pp_1_3_2;
  wire pp_1_3_3;
  wire pp_1_4_0;
  wire pp_1_4_1;
  wire pp_1_4_2;
  wire pp_1_5_0;
  wire pp_1_5_1;
  wire pp_1_5_2;
  wire pp_1_6_0;
  wire pp_1_6_1;
  wire pp_1_6_2;
  wire pp_1_6_3;
  wire pp_1_6_4;
  wire pp_1_6_5;
  wire pp_1_6_6;
  wire pp_1_6_7;
  wire pp_1_6_8;
  wire pp_1_7_0;
  wire pp_1_7_1;
  wire pp_1_7_2;
  wire pp_1_8_0;
  wire pp_1_8_1;
  wire pp_1_8_2;
  wire pp_1_8_3;
  wire pp_1_8_4;
  wire pp_1_8_5;
  wire pp_1_8_6;
  wire pp_1_8_7;
  wire pp_1_8_8;
  wire pp_1_8_9;
  wire pp_1_8_10;
  wire pp_1_8_11;
  wire pp_1_9_0;
  wire pp_1_9_1;
  wire pp_1_9_2;
  wire pp_1_9_3;
  wire pp_1_9_4;
  wire pp_1_9_5;
  wire pp_1_9_6;
  wire pp_1_9_7;
  wire pp_1_9_8;
  wire pp_1_9_9;
  wire pp_1_10_0;
  wire pp_1_10_1;
  wire pp_1_10_2;
  wire pp_1_10_3;
  wire pp_1_10_4;
  wire pp_1_11_0;
  wire pp_1_11_1;
  wire pp_1_11_2;
  wire pp_1_11_3;
  wire pp_1_11_4;
  wire pp_1_11_5;
  wire pp_1_11_6;
  wire pp_1_11_7;
  wire pp_1_11_8;
  wire pp_1_12_0;
  wire pp_1_12_1;
  wire pp_1_12_2;
  wire pp_1_12_3;
  wire pp_1_12_4;
  wire pp_1_12_5;
  wire pp_1_12_6;
  wire pp_1_12_7;
  wire pp_1_12_8;
  wire pp_1_13_0;
  wire pp_1_13_1;
  wire pp_1_13_2;
  wire pp_1_13_3;
  wire pp_1_13_4;
  wire pp_1_13_5;
  wire pp_1_13_6;
  wire pp_1_13_7;
  wire pp_1_13_8;
  wire pp_1_14_0;
  wire pp_1_14_1;
  wire pp_1_14_2;
  wire pp_1_14_3;
  wire pp_1_14_4;
  wire pp_1_14_5;
  wire pp_1_14_6;
  wire pp_1_14_7;
  wire pp_1_14_8;
  wire pp_1_14_9;
  wire pp_1_14_10;
  wire pp_1_14_11;
  wire pp_1_14_12;
  wire pp_1_14_13;
  wire pp_1_14_14;
  wire pp_1_14_15;
  wire pp_1_14_16;
  wire pp_1_14_17;
  wire pp_1_14_18;
  wire pp_1_14_19;
  wire pp_1_15_0;
  wire pp_1_15_1;
  wire pp_1_15_2;
  wire pp_1_15_3;
  wire pp_1_15_4;
  wire pp_1_15_5;
  wire pp_1_16_0;
  wire pp_1_16_1;
  wire pp_1_16_2;
  wire pp_1_16_3;
  wire pp_1_16_4;
  wire pp_1_16_5;
  wire pp_1_16_6;
  wire pp_1_16_7;
  wire pp_1_16_8;
  wire pp_1_16_9;
  wire pp_1_16_10;
  wire pp_1_16_11;
  wire pp_1_16_12;
  wire pp_1_16_13;
  wire pp_1_16_14;
  wire pp_1_16_15;
  wire pp_1_16_16;
  wire pp_1_16_17;
  wire pp_1_16_18;
  wire pp_1_16_19;
  wire pp_1_16_20;
  wire pp_1_17_0;
  wire pp_1_17_1;
  wire pp_1_17_2;
  wire pp_1_17_3;
  wire pp_1_17_4;
  wire pp_1_17_5;
  wire pp_1_18_0;
  wire pp_1_18_1;
  wire pp_1_18_2;
  wire pp_1_18_3;
  wire pp_1_18_4;
  wire pp_1_18_5;
  wire pp_1_18_6;
  wire pp_1_18_7;
  wire pp_1_18_8;
  wire pp_1_19_0;
  wire pp_1_19_1;
  wire pp_1_19_2;
  wire pp_1_19_3;
  wire pp_1_19_4;
  wire pp_1_19_5;
  wire pp_1_19_6;
  wire pp_1_19_7;
  wire pp_1_20_0;
  wire pp_1_20_1;
  wire pp_1_20_2;
  wire pp_1_20_3;
  wire pp_1_20_4;
  wire pp_1_20_5;
  wire pp_1_20_6;
  wire pp_1_20_7;
  wire pp_1_20_8;
  wire pp_1_21_0;
  wire pp_1_21_1;
  wire pp_1_21_2;
  wire pp_1_21_3;
  wire pp_1_21_4;
  wire pp_1_21_5;
  wire pp_1_21_6;
  wire pp_1_22_0;
  wire pp_1_22_1;
  wire pp_1_22_2;
  wire pp_1_22_3;
  wire pp_1_22_4;
  wire pp_1_22_5;
  wire pp_1_23_0;
  wire pp_1_23_1;
  wire pp_1_23_2;
  wire pp_1_23_3;
  wire pp_1_23_4;
  wire pp_1_23_5;
  wire pp_1_23_6;
  wire pp_1_23_7;
  wire pp_1_23_8;
  wire pp_1_23_9;
  wire pp_1_23_10;
  wire pp_1_24_0;
  wire pp_1_24_1;
  wire pp_1_24_2;
  wire pp_1_24_3;
  wire pp_1_24_4;
  wire pp_1_25_0;
  wire pp_1_25_1;
  wire pp_1_25_2;
  wire pp_1_26_0;
  wire pp_1_26_1;
  wire pp_1_26_2;
  wire pp_1_26_3;
  wire pp_1_26_4;
  wire pp_1_26_5;
  wire pp_1_26_6;
  wire pp_1_27_0;
  wire pp_1_27_1;
  wire pp_1_27_2;
  wire pp_1_27_3;
  wire pp_1_28_0;
  wire pp_1_29_0;
  wire pp_1_29_1;
  wire pp_1_29_2;
  wire pp_1_30_0;
  wire pp_1_31_0;
  wire pp_2_0_0;
  wire pp_2_1_0;
  wire pp_2_1_1;
  wire pp_2_2_0;
  wire pp_2_2_1;
  wire pp_2_2_2;
  wire pp_2_3_0;
  wire pp_2_3_1;
  wire pp_2_4_0;
  wire pp_2_4_1;
  wire pp_2_5_0;
  wire pp_2_5_1;
  wire pp_2_6_0;
  wire pp_2_6_1;
  wire pp_2_6_2;
  wire pp_2_6_3;
  wire pp_2_7_0;
  wire pp_2_7_1;
  wire pp_2_7_2;
  wire pp_2_7_3;
  wire pp_2_8_0;
  wire pp_2_8_1;
  wire pp_2_8_2;
  wire pp_2_8_3;
  wire pp_2_8_4;
  wire pp_2_9_0;
  wire pp_2_9_1;
  wire pp_2_9_2;
  wire pp_2_9_3;
  wire pp_2_9_4;
  wire pp_2_9_5;
  wire pp_2_9_6;
  wire pp_2_9_7;
  wire pp_2_10_0;
  wire pp_2_10_1;
  wire pp_2_10_2;
  wire pp_2_10_3;
  wire pp_2_10_4;
  wire pp_2_10_5;
  wire pp_2_11_0;
  wire pp_2_11_1;
  wire pp_2_11_2;
  wire pp_2_11_3;
  wire pp_2_12_0;
  wire pp_2_12_1;
  wire pp_2_12_2;
  wire pp_2_12_3;
  wire pp_2_12_4;
  wire pp_2_12_5;
  wire pp_2_13_0;
  wire pp_2_13_1;
  wire pp_2_13_2;
  wire pp_2_13_3;
  wire pp_2_13_4;
  wire pp_2_13_5;
  wire pp_2_14_0;
  wire pp_2_14_1;
  wire pp_2_14_2;
  wire pp_2_14_3;
  wire pp_2_14_4;
  wire pp_2_14_5;
  wire pp_2_14_6;
  wire pp_2_14_7;
  wire pp_2_14_8;
  wire pp_2_14_9;
  wire pp_2_15_0;
  wire pp_2_15_1;
  wire pp_2_15_2;
  wire pp_2_15_3;
  wire pp_2_15_4;
  wire pp_2_15_5;
  wire pp_2_15_6;
  wire pp_2_15_7;
  wire pp_2_15_8;
  wire pp_2_16_0;
  wire pp_2_16_1;
  wire pp_2_16_2;
  wire pp_2_16_3;
  wire pp_2_16_4;
  wire pp_2_16_5;
  wire pp_2_16_6;
  wire pp_2_16_7;
  wire pp_2_16_8;
  wire pp_2_17_0;
  wire pp_2_17_1;
  wire pp_2_17_2;
  wire pp_2_17_3;
  wire pp_2_17_4;
  wire pp_2_17_5;
  wire pp_2_17_6;
  wire pp_2_17_7;
  wire pp_2_17_8;
  wire pp_2_18_0;
  wire pp_2_18_1;
  wire pp_2_18_2;
  wire pp_2_18_3;
  wire pp_2_18_4;
  wire pp_2_19_0;
  wire pp_2_19_1;
  wire pp_2_19_2;
  wire pp_2_19_3;
  wire pp_2_19_4;
  wire pp_2_19_5;
  wire pp_2_19_6;
  wire pp_2_20_0;
  wire pp_2_20_1;
  wire pp_2_20_2;
  wire pp_2_20_3;
  wire pp_2_20_4;
  wire pp_2_21_0;
  wire pp_2_21_1;
  wire pp_2_21_2;
  wire pp_2_21_3;
  wire pp_2_21_4;
  wire pp_2_21_5;
  wire pp_2_22_0;
  wire pp_2_22_1;
  wire pp_2_22_2;
  wire pp_2_22_3;
  wire pp_2_23_0;
  wire pp_2_23_1;
  wire pp_2_23_2;
  wire pp_2_23_3;
  wire pp_2_23_4;
  wire pp_2_23_5;
  wire pp_2_23_6;
  wire pp_2_24_0;
  wire pp_2_24_1;
  wire pp_2_24_2;
  wire pp_2_24_3;
  wire pp_2_24_4;
  wire pp_2_24_5;
  wire pp_2_25_0;
  wire pp_2_25_1;
  wire pp_2_26_0;
  wire pp_2_26_1;
  wire pp_2_26_2;
  wire pp_2_26_3;
  wire pp_2_27_0;
  wire pp_2_27_1;
  wire pp_2_27_2;
  wire pp_2_27_3;
  wire pp_2_28_0;
  wire pp_2_28_1;
  wire pp_2_29_0;
  wire pp_2_30_0;
  wire pp_2_30_1;
  wire pp_2_31_0;
  wire pp_3_0_0;
  wire pp_3_1_0;
  wire pp_3_1_1;
  wire pp_3_2_0;
  wire pp_3_2_1;
  wire pp_3_2_2;
  wire pp_3_3_0;
  wire pp_3_3_1;
  wire pp_3_4_0;
  wire pp_3_4_1;
  wire pp_3_5_0;
  wire pp_3_5_1;
  wire pp_3_6_0;
  wire pp_3_6_1;
  wire pp_3_6_2;
  wire pp_3_6_3;
  wire pp_3_7_0;
  wire pp_3_7_1;
  wire pp_3_8_0;
  wire pp_3_8_1;
  wire pp_3_8_2;
  wire pp_3_8_3;
  wire pp_3_8_4;
  wire pp_3_8_5;
  wire pp_3_9_0;
  wire pp_3_9_1;
  wire pp_3_9_2;
  wire pp_3_10_0;
  wire pp_3_10_1;
  wire pp_3_10_2;
  wire pp_3_10_3;
  wire pp_3_10_4;
  wire pp_3_11_0;
  wire pp_3_11_1;
  wire pp_3_11_2;
  wire pp_3_11_3;
  wire pp_3_12_0;
  wire pp_3_12_1;
  wire pp_3_12_2;
  wire pp_3_13_0;
  wire pp_3_13_1;
  wire pp_3_13_2;
  wire pp_3_13_3;
  wire pp_3_14_0;
  wire pp_3_14_1;
  wire pp_3_14_2;
  wire pp_3_14_3;
  wire pp_3_14_4;
  wire pp_3_14_5;
  wire pp_3_15_0;
  wire pp_3_15_1;
  wire pp_3_15_2;
  wire pp_3_15_3;
  wire pp_3_15_4;
  wire pp_3_15_5;
  wire pp_3_16_0;
  wire pp_3_16_1;
  wire pp_3_16_2;
  wire pp_3_16_3;
  wire pp_3_16_4;
  wire pp_3_16_5;
  wire pp_3_17_0;
  wire pp_3_17_1;
  wire pp_3_17_2;
  wire pp_3_17_3;
  wire pp_3_17_4;
  wire pp_3_17_5;
  wire pp_3_18_0;
  wire pp_3_18_1;
  wire pp_3_18_2;
  wire pp_3_18_3;
  wire pp_3_18_4;
  wire pp_3_18_5;
  wire pp_3_19_0;
  wire pp_3_19_1;
  wire pp_3_19_2;
  wire pp_3_19_3;
  wire pp_3_19_4;
  wire pp_3_19_5;
  wire pp_3_20_0;
  wire pp_3_20_1;
  wire pp_3_20_2;
  wire pp_3_20_3;
  wire pp_3_21_0;
  wire pp_3_21_1;
  wire pp_3_21_2;
  wire pp_3_22_0;
  wire pp_3_22_1;
  wire pp_3_22_2;
  wire pp_3_22_3;
  wire pp_3_22_4;
  wire pp_3_22_5;
  wire pp_3_23_0;
  wire pp_3_23_1;
  wire pp_3_23_2;
  wire pp_3_24_0;
  wire pp_3_24_1;
  wire pp_3_24_2;
  wire pp_3_24_3;
  wire pp_3_24_4;
  wire pp_3_24_5;
  wire pp_3_25_0;
  wire pp_3_25_1;
  wire pp_3_25_2;
  wire pp_3_26_0;
  wire pp_3_26_1;
  wire pp_3_26_2;
  wire pp_3_26_3;
  wire pp_3_27_0;
  wire pp_3_27_1;
  wire pp_3_28_0;
  wire pp_3_28_1;
  wire pp_3_28_2;
  wire pp_3_29_0;
  wire pp_3_30_0;
  wire pp_3_30_1;
  wire pp_3_31_0;
  wire pp_4_0_0;
  wire pp_4_1_0;
  wire pp_4_1_1;
  wire pp_4_2_0;
  wire pp_4_2_1;
  wire pp_4_2_2;
  wire pp_4_3_0;
  wire pp_4_3_1;
  wire pp_4_4_0;
  wire pp_4_4_1;
  wire pp_4_5_0;
  wire pp_4_5_1;
  wire pp_4_6_0;
  wire pp_4_6_1;
  wire pp_4_7_0;
  wire pp_4_7_1;
  wire pp_4_7_2;
  wire pp_4_8_0;
  wire pp_4_8_1;
  wire pp_4_9_0;
  wire pp_4_9_1;
  wire pp_4_9_2;
  wire pp_4_10_0;
  wire pp_4_10_1;
  wire pp_4_10_2;
  wire pp_4_11_0;
  wire pp_4_11_1;
  wire pp_4_11_2;
  wire pp_4_11_3;
  wire pp_4_11_4;
  wire pp_4_11_5;
  wire pp_4_12_0;
  wire pp_4_12_1;
  wire pp_4_12_2;
  wire pp_4_13_0;
  wire pp_4_13_1;
  wire pp_4_13_2;
  wire pp_4_13_3;
  wire pp_4_14_0;
  wire pp_4_14_1;
  wire pp_4_15_0;
  wire pp_4_15_1;
  wire pp_4_15_2;
  wire pp_4_15_3;
  wire pp_4_15_4;
  wire pp_4_15_5;
  wire pp_4_16_0;
  wire pp_4_16_1;
  wire pp_4_16_2;
  wire pp_4_17_0;
  wire pp_4_17_1;
  wire pp_4_17_2;
  wire pp_4_17_3;
  wire pp_4_18_0;
  wire pp_4_18_1;
  wire pp_4_18_2;
  wire pp_4_18_3;
  wire pp_4_19_0;
  wire pp_4_19_1;
  wire pp_4_19_2;
  wire pp_4_19_3;
  wire pp_4_20_0;
  wire pp_4_20_1;
  wire pp_4_20_2;
  wire pp_4_20_3;
  wire pp_4_20_4;
  wire pp_4_20_5;
  wire pp_4_21_0;
  wire pp_4_22_0;
  wire pp_4_22_1;
  wire pp_4_22_2;
  wire pp_4_23_0;
  wire pp_4_23_1;
  wire pp_4_23_2;
  wire pp_4_23_3;
  wire pp_4_23_4;
  wire pp_4_24_0;
  wire pp_4_24_1;
  wire pp_4_25_0;
  wire pp_4_25_1;
  wire pp_4_25_2;
  wire pp_4_26_0;
  wire pp_4_26_1;
  wire pp_4_26_2;
  wire pp_4_27_0;
  wire pp_4_27_1;
  wire pp_4_27_2;
  wire pp_4_28_0;
  wire pp_4_28_1;
  wire pp_4_28_2;
  wire pp_4_29_0;
  wire pp_4_30_0;
  wire pp_4_30_1;
  wire pp_4_31_0;
  wire pp_5_0_0;
  wire pp_5_1_0;
  wire pp_5_1_1;
  wire pp_5_2_0;
  wire pp_5_2_1;
  wire pp_5_2_2;
  wire pp_5_3_0;
  wire pp_5_4_0;
  wire pp_5_4_1;
  wire pp_5_5_0;
  wire pp_5_5_1;
  wire pp_5_6_0;
  wire pp_5_6_1;
  wire pp_5_7_0;
  wire pp_5_7_1;
  wire pp_5_8_0;
  wire pp_5_8_1;
  wire pp_5_8_2;
  wire pp_5_9_0;
  wire pp_5_9_1;
  wire pp_5_9_2;
  wire pp_5_10_0;
  wire pp_5_11_0;
  wire pp_5_11_1;
  wire pp_5_11_2;
  wire pp_5_12_0;
  wire pp_5_12_1;
  wire pp_5_12_2;
  wire pp_5_13_0;
  wire pp_5_13_1;
  wire pp_5_13_2;
  wire pp_5_14_0;
  wire pp_5_14_1;
  wire pp_5_14_2;
  wire pp_5_15_0;
  wire pp_5_15_1;
  wire pp_5_16_0;
  wire pp_5_16_1;
  wire pp_5_16_2;
  wire pp_5_17_0;
  wire pp_5_17_1;
  wire pp_5_17_2;
  wire pp_5_18_0;
  wire pp_5_18_1;
  wire pp_5_18_2;
  wire pp_5_19_0;
  wire pp_5_19_1;
  wire pp_5_19_2;
  wire pp_5_20_0;
  wire pp_5_20_1;
  wire pp_5_20_2;
  wire pp_5_21_0;
  wire pp_5_21_1;
  wire pp_5_21_2;
  wire pp_5_22_0;
  wire pp_5_22_1;
  wire pp_5_22_2;
  wire pp_5_23_0;
  wire pp_5_23_1;
  wire pp_5_23_2;
  wire pp_5_24_0;
  wire pp_5_24_1;
  wire pp_5_24_2;
  wire pp_5_25_0;
  wire pp_5_26_0;
  wire pp_5_26_1;
  wire pp_5_26_2;
  wire pp_5_26_3;
  wire pp_5_27_0;
  wire pp_5_28_0;
  wire pp_5_28_1;
  wire pp_5_28_2;
  wire pp_5_28_3;
  wire pp_5_29_0;
  wire pp_5_30_0;
  wire pp_5_30_1;
  wire pp_5_31_0;
  wire pp_6_0_0;
  wire pp_6_1_0;
  wire pp_6_1_1;
  wire pp_6_2_0;
  wire pp_6_2_1;
  wire pp_6_3_0;
  wire pp_6_3_1;
  wire pp_6_4_0;
  wire pp_6_4_1;
  wire pp_6_5_0;
  wire pp_6_5_1;
  wire pp_6_6_0;
  wire pp_6_6_1;
  wire pp_6_7_0;
  wire pp_6_7_1;
  wire pp_6_8_0;
  wire pp_6_8_1;
  wire pp_6_9_0;
  wire pp_6_9_1;
  wire pp_6_10_0;
  wire pp_6_10_1;
  wire pp_6_11_0;
  wire pp_6_11_1;
  wire pp_6_12_0;
  wire pp_6_12_1;
  wire pp_6_13_0;
  wire pp_6_13_1;
  wire pp_6_14_0;
  wire pp_6_14_1;
  wire pp_6_15_0;
  wire pp_6_15_1;
  wire pp_6_16_0;
  wire pp_6_16_1;
  wire pp_6_17_0;
  wire pp_6_17_1;
  wire pp_6_18_0;
  wire pp_6_18_1;
  wire pp_6_19_0;
  wire pp_6_19_1;
  wire pp_6_20_0;
  wire pp_6_20_1;
  wire pp_6_21_0;
  wire pp_6_21_1;
  wire pp_6_22_0;
  wire pp_6_22_1;
  wire pp_6_23_0;
  wire pp_6_23_1;
  wire pp_6_24_0;
  wire pp_6_24_1;
  wire pp_6_25_0;
  wire pp_6_25_1;
  wire pp_6_26_0;
  wire pp_6_26_1;
  wire pp_6_27_0;
  wire pp_6_27_1;
  wire pp_6_28_0;
  wire pp_6_28_1;
  wire pp_6_29_0;
  wire pp_6_29_1;
  wire pp_6_30_0;
  wire pp_6_30_1;
  wire pp_6_31_0;
  assign pp_0_0_0 = pp_0_0;
  assign pp_0_1_0 = pp_0_1;
  assign pp_0_1_1 = pp_1_1;
  assign pp_0_2_0 = pp_0_2;
  assign pp_0_2_1 = pp_1_2;
  assign pp_0_2_2 = pp_2_2;
  assign pp_0_3_0 = pp_0_3;
  assign pp_0_3_1 = pp_1_3;
  assign pp_0_3_2 = pp_2_3;
  assign pp_0_3_3 = pp_3_3;
  assign pp_0_4_0 = pp_0_4;
  assign pp_0_4_1 = pp_1_4;
  assign pp_0_4_2 = pp_2_4;
  assign pp_0_4_3 = pp_3_4;
  assign pp_0_4_4 = pp_4_4;
  assign pp_0_5_0 = pp_0_5;
  assign pp_0_5_1 = pp_1_5;
  assign pp_0_5_2 = pp_2_5;
  assign pp_0_5_3 = pp_3_5;
  assign pp_0_5_4 = pp_4_5;
  assign pp_0_5_5 = pp_5_5;
  assign pp_0_6_0 = pp_0_6;
  assign pp_0_6_1 = pp_1_6;
  assign pp_0_6_2 = pp_2_6;
  assign pp_0_6_3 = pp_3_6;
  assign pp_0_6_4 = pp_4_6;
  assign pp_0_6_5 = pp_5_6;
  assign pp_0_6_6 = pp_6_6;
  assign pp_0_7_0 = pp_0_7;
  assign pp_0_7_1 = pp_1_7;
  assign pp_0_7_2 = pp_2_7;
  assign pp_0_7_3 = pp_3_7;
  assign pp_0_7_4 = pp_4_7;
  assign pp_0_7_5 = pp_5_7;
  assign pp_0_7_6 = pp_6_7;
  assign pp_0_7_7 = pp_7_7;
  assign pp_0_8_0 = pp_0_8;
  assign pp_0_8_1 = pp_1_8;
  assign pp_0_8_2 = pp_2_8;
  assign pp_0_8_3 = pp_3_8;
  assign pp_0_8_4 = pp_4_8;
  assign pp_0_8_5 = pp_5_8;
  assign pp_0_8_6 = pp_6_8;
  assign pp_0_8_7 = pp_7_8;
  assign pp_0_8_8 = pp_8_8;
  assign pp_0_9_0 = pp_0_9;
  assign pp_0_9_1 = pp_1_9;
  assign pp_0_9_2 = pp_2_9;
  assign pp_0_9_3 = pp_3_9;
  assign pp_0_9_4 = pp_4_9;
  assign pp_0_9_5 = pp_5_9;
  assign pp_0_9_6 = pp_6_9;
  assign pp_0_9_7 = pp_7_9;
  assign pp_0_9_8 = pp_8_9;
  assign pp_0_9_9 = pp_9_9;
  assign pp_0_10_0 = pp_0_10;
  assign pp_0_10_1 = pp_1_10;
  assign pp_0_10_2 = pp_2_10;
  assign pp_0_10_3 = pp_3_10;
  assign pp_0_10_4 = pp_4_10;
  assign pp_0_10_5 = pp_5_10;
  assign pp_0_10_6 = pp_6_10;
  assign pp_0_10_7 = pp_7_10;
  assign pp_0_10_8 = pp_8_10;
  assign pp_0_10_9 = pp_9_10;
  assign pp_0_10_10 = pp_10_10;
  assign pp_0_11_0 = pp_0_11;
  assign pp_0_11_1 = pp_1_11;
  assign pp_0_11_2 = pp_2_11;
  assign pp_0_11_3 = pp_3_11;
  assign pp_0_11_4 = pp_4_11;
  assign pp_0_11_5 = pp_5_11;
  assign pp_0_11_6 = pp_6_11;
  assign pp_0_11_7 = pp_7_11;
  assign pp_0_11_8 = pp_8_11;
  assign pp_0_11_9 = pp_9_11;
  assign pp_0_11_10 = pp_10_11;
  assign pp_0_11_11 = pp_11_11;
  assign pp_0_12_0 = pp_0_12;
  assign pp_0_12_1 = pp_1_12;
  assign pp_0_12_2 = pp_2_12;
  assign pp_0_12_3 = pp_3_12;
  assign pp_0_12_4 = pp_4_12;
  assign pp_0_12_5 = pp_5_12;
  assign pp_0_12_6 = pp_6_12;
  assign pp_0_12_7 = pp_7_12;
  assign pp_0_12_8 = pp_8_12;
  assign pp_0_12_9 = pp_9_12;
  assign pp_0_12_10 = pp_10_12;
  assign pp_0_12_11 = pp_11_12;
  assign pp_0_12_12 = pp_12_12;
  assign pp_0_13_0 = pp_0_13;
  assign pp_0_13_1 = pp_1_13;
  assign pp_0_13_2 = pp_2_13;
  assign pp_0_13_3 = pp_3_13;
  assign pp_0_13_4 = pp_4_13;
  assign pp_0_13_5 = pp_5_13;
  assign pp_0_13_6 = pp_6_13;
  assign pp_0_13_7 = pp_7_13;
  assign pp_0_13_8 = pp_8_13;
  assign pp_0_13_9 = pp_9_13;
  assign pp_0_13_10 = pp_10_13;
  assign pp_0_13_11 = pp_11_13;
  assign pp_0_13_12 = pp_12_13;
  assign pp_0_13_13 = pp_13_13;
  assign pp_0_14_0 = pp_0_14;
  assign pp_0_14_1 = pp_1_14;
  assign pp_0_14_2 = pp_2_14;
  assign pp_0_14_3 = pp_3_14;
  assign pp_0_14_4 = pp_4_14;
  assign pp_0_14_5 = pp_5_14;
  assign pp_0_14_6 = pp_6_14;
  assign pp_0_14_7 = pp_7_14;
  assign pp_0_14_8 = pp_8_14;
  assign pp_0_14_9 = pp_9_14;
  assign pp_0_14_10 = pp_10_14;
  assign pp_0_14_11 = pp_11_14;
  assign pp_0_14_12 = pp_12_14;
  assign pp_0_14_13 = pp_13_14;
  assign pp_0_14_14 = pp_14_14;
  assign pp_0_15_0 = pp_0_15;
  assign pp_0_15_1 = pp_1_15;
  assign pp_0_15_2 = pp_2_15;
  assign pp_0_15_3 = pp_3_15;
  assign pp_0_15_4 = pp_4_15;
  assign pp_0_15_5 = pp_5_15;
  assign pp_0_15_6 = pp_6_15;
  assign pp_0_15_7 = pp_7_15;
  assign pp_0_15_8 = pp_8_15;
  assign pp_0_15_9 = pp_9_15;
  assign pp_0_15_10 = pp_10_15;
  assign pp_0_15_11 = pp_11_15;
  assign pp_0_15_12 = pp_12_15;
  assign pp_0_15_13 = pp_13_15;
  assign pp_0_15_14 = pp_14_15;
  assign pp_0_15_15 = pp_15_15;
  assign pp_0_16_0 = pp_0_16;
  assign pp_0_16_1 = pp_1_16;
  assign pp_0_16_2 = pp_2_16;
  assign pp_0_16_3 = pp_3_16;
  assign pp_0_16_4 = pp_4_16;
  assign pp_0_16_5 = pp_5_16;
  assign pp_0_16_6 = pp_6_16;
  assign pp_0_16_7 = pp_7_16;
  assign pp_0_16_8 = pp_8_16;
  assign pp_0_16_9 = pp_9_16;
  assign pp_0_16_10 = pp_10_16;
  assign pp_0_16_11 = pp_11_16;
  assign pp_0_16_12 = pp_12_16;
  assign pp_0_16_13 = pp_13_16;
  assign pp_0_16_14 = pp_14_16;
  assign pp_0_16_15 = pp_15_16;
  assign pp_0_17_0 = pp_2_17;
  assign pp_0_17_1 = pp_3_17;
  assign pp_0_17_2 = pp_4_17;
  assign pp_0_17_3 = pp_5_17;
  assign pp_0_17_4 = pp_6_17;
  assign pp_0_17_5 = pp_7_17;
  assign pp_0_17_6 = pp_8_17;
  assign pp_0_17_7 = pp_9_17;
  assign pp_0_17_8 = pp_10_17;
  assign pp_0_17_9 = pp_11_17;
  assign pp_0_17_10 = pp_12_17;
  assign pp_0_17_11 = pp_13_17;
  assign pp_0_17_12 = pp_14_17;
  assign pp_0_17_13 = pp_15_17;
  assign pp_0_18_0 = pp_3_18;
  assign pp_0_18_1 = pp_4_18;
  assign pp_0_18_2 = pp_5_18;
  assign pp_0_18_3 = pp_6_18;
  assign pp_0_18_4 = pp_7_18;
  assign pp_0_18_5 = pp_8_18;
  assign pp_0_18_6 = pp_9_18;
  assign pp_0_18_7 = pp_10_18;
  assign pp_0_18_8 = pp_11_18;
  assign pp_0_18_9 = pp_12_18;
  assign pp_0_18_10 = pp_13_18;
  assign pp_0_18_11 = pp_14_18;
  assign pp_0_18_12 = pp_15_18;
  assign pp_0_19_0 = pp_4_19;
  assign pp_0_19_1 = pp_5_19;
  assign pp_0_19_2 = pp_6_19;
  assign pp_0_19_3 = pp_7_19;
  assign pp_0_19_4 = pp_8_19;
  assign pp_0_19_5 = pp_9_19;
  assign pp_0_19_6 = pp_10_19;
  assign pp_0_19_7 = pp_11_19;
  assign pp_0_19_8 = pp_12_19;
  assign pp_0_19_9 = pp_13_19;
  assign pp_0_19_10 = pp_14_19;
  assign pp_0_19_11 = pp_15_19;
  assign pp_0_20_0 = pp_5_20;
  assign pp_0_20_1 = pp_6_20;
  assign pp_0_20_2 = pp_7_20;
  assign pp_0_20_3 = pp_8_20;
  assign pp_0_20_4 = pp_9_20;
  assign pp_0_20_5 = pp_10_20;
  assign pp_0_20_6 = pp_11_20;
  assign pp_0_20_7 = pp_12_20;
  assign pp_0_20_8 = pp_13_20;
  assign pp_0_20_9 = pp_14_20;
  assign pp_0_20_10 = pp_15_20;
  assign pp_0_21_0 = pp_6_21;
  assign pp_0_21_1 = pp_7_21;
  assign pp_0_21_2 = pp_8_21;
  assign pp_0_21_3 = pp_9_21;
  assign pp_0_21_4 = pp_10_21;
  assign pp_0_21_5 = pp_11_21;
  assign pp_0_21_6 = pp_12_21;
  assign pp_0_21_7 = pp_13_21;
  assign pp_0_21_8 = pp_14_21;
  assign pp_0_21_9 = pp_15_21;
  assign pp_0_22_0 = pp_7_22;
  assign pp_0_22_1 = pp_8_22;
  assign pp_0_22_2 = pp_9_22;
  assign pp_0_22_3 = pp_10_22;
  assign pp_0_22_4 = pp_11_22;
  assign pp_0_22_5 = pp_12_22;
  assign pp_0_22_6 = pp_13_22;
  assign pp_0_22_7 = pp_14_22;
  assign pp_0_22_8 = pp_15_22;
  assign pp_0_23_0 = pp_8_23;
  assign pp_0_23_1 = pp_9_23;
  assign pp_0_23_2 = pp_10_23;
  assign pp_0_23_3 = pp_11_23;
  assign pp_0_23_4 = pp_12_23;
  assign pp_0_23_5 = pp_13_23;
  assign pp_0_23_6 = pp_14_23;
  assign pp_0_23_7 = pp_15_23;
  assign pp_0_24_0 = pp_9_24;
  assign pp_0_24_1 = pp_10_24;
  assign pp_0_24_2 = pp_11_24;
  assign pp_0_24_3 = pp_12_24;
  assign pp_0_24_4 = pp_13_24;
  assign pp_0_24_5 = pp_14_24;
  assign pp_0_24_6 = pp_15_24;
  assign pp_0_25_0 = pp_10_25;
  assign pp_0_25_1 = pp_11_25;
  assign pp_0_25_2 = pp_12_25;
  assign pp_0_25_3 = pp_13_25;
  assign pp_0_25_4 = pp_14_25;
  assign pp_0_25_5 = pp_15_25;
  assign pp_0_26_0 = pp_11_26;
  assign pp_0_26_1 = pp_12_26;
  assign pp_0_26_2 = pp_13_26;
  assign pp_0_26_3 = pp_14_26;
  assign pp_0_26_4 = pp_15_26;
  assign pp_0_27_0 = pp_12_27;
  assign pp_0_27_1 = pp_13_27;
  assign pp_0_27_2 = pp_14_27;
  assign pp_0_27_3 = pp_15_27;
  assign pp_0_28_0 = pp_13_28;
  assign pp_0_28_1 = pp_14_28;
  assign pp_0_28_2 = pp_15_28;
  assign pp_0_29_0 = pp_14_29;
  assign pp_0_29_1 = pp_15_29;
  assign pp_0_30_0 = pp_15_30;
  assign pp_0_31_0 = pp_15_31;

  assign pp_1_0_0 = pp_0_0_0;
  assign pp_1_1_0 = pp_0_1_0;
  assign pp_1_1_1 = pp_0_1_1;
  assign pp_1_2_0 = pp_0_2_0;
  assign pp_1_2_1 = pp_0_2_1;
  assign pp_1_2_2 = pp_0_2_2;
  assign pp_1_3_0 = pp_0_3_0;
  assign pp_1_3_1 = pp_0_3_1;
  assign pp_1_3_2 = pp_0_3_2;
  assign pp_1_3_3 = pp_0_3_3;
  MG_FA fa_0_4_0(
    .a(pp_0_4_0),
    .b(pp_0_4_1),
    .cin(pp_0_4_2),
    .sum(pp_1_4_0),
    .cout(pp_1_5_0)
  );

  assign pp_1_4_1 = pp_0_4_3;
  assign pp_1_4_2 = pp_0_4_4;
  MG_FA fa_0_5_0(
    .a(pp_0_5_0),
    .b(pp_0_5_1),
    .cin(pp_0_5_2),
    .sum(pp_1_5_1),
    .cout(pp_1_6_0)
  );

  MG_FA fa_0_5_1(
    .a(pp_0_5_3),
    .b(pp_0_5_4),
    .cin(pp_0_5_5),
    .sum(pp_1_5_2),
    .cout(pp_1_6_1)
  );

  assign pp_1_6_2 = pp_0_6_0;
  assign pp_1_6_3 = pp_0_6_1;
  assign pp_1_6_4 = pp_0_6_2;
  assign pp_1_6_5 = pp_0_6_3;
  assign pp_1_6_6 = pp_0_6_4;
  assign pp_1_6_7 = pp_0_6_5;
  assign pp_1_6_8 = pp_0_6_6;
  MG_FA fa_0_7_0(
    .a(pp_0_7_0),
    .b(pp_0_7_1),
    .cin(pp_0_7_2),
    .sum(pp_1_7_0),
    .cout(pp_1_8_0)
  );

  MG_FA fa_0_7_1(
    .a(pp_0_7_3),
    .b(pp_0_7_4),
    .cin(pp_0_7_5),
    .sum(pp_1_7_1),
    .cout(pp_1_8_1)
  );

  MG_HA ha_0_7_2(
    .a(pp_0_7_6),
    .b(pp_0_7_7),
    .sum(pp_1_7_2),
    .cout(pp_1_8_2)
  );

  assign pp_1_8_3 = pp_0_8_0;
  assign pp_1_8_4 = pp_0_8_1;
  assign pp_1_8_5 = pp_0_8_2;
  assign pp_1_8_6 = pp_0_8_3;
  assign pp_1_8_7 = pp_0_8_4;
  assign pp_1_8_8 = pp_0_8_5;
  assign pp_1_8_9 = pp_0_8_6;
  assign pp_1_8_10 = pp_0_8_7;
  assign pp_1_8_11 = pp_0_8_8;
  assign pp_1_9_0 = pp_0_9_0;
  assign pp_1_9_1 = pp_0_9_1;
  assign pp_1_9_2 = pp_0_9_2;
  assign pp_1_9_3 = pp_0_9_3;
  assign pp_1_9_4 = pp_0_9_4;
  assign pp_1_9_5 = pp_0_9_5;
  assign pp_1_9_6 = pp_0_9_6;
  assign pp_1_9_7 = pp_0_9_7;
  assign pp_1_9_8 = pp_0_9_8;
  assign pp_1_9_9 = pp_0_9_9;
  MG_FA fa_0_10_0(
    .a(pp_0_10_0),
    .b(pp_0_10_1),
    .cin(pp_0_10_2),
    .sum(pp_1_10_0),
    .cout(pp_1_11_0)
  );

  MG_FA fa_0_10_1(
    .a(pp_0_10_3),
    .b(pp_0_10_4),
    .cin(pp_0_10_5),
    .sum(pp_1_10_1),
    .cout(pp_1_11_1)
  );

  MG_FA fa_0_10_2(
    .a(pp_0_10_6),
    .b(pp_0_10_7),
    .cin(pp_0_10_8),
    .sum(pp_1_10_2),
    .cout(pp_1_11_2)
  );

  assign pp_1_10_3 = pp_0_10_9;
  assign pp_1_10_4 = pp_0_10_10;
  MG_FA fa_0_11_0(
    .a(pp_0_11_0),
    .b(pp_0_11_1),
    .cin(pp_0_11_2),
    .sum(pp_1_11_3),
    .cout(pp_1_12_0)
  );

  MG_FA fa_0_11_1(
    .a(pp_0_11_3),
    .b(pp_0_11_4),
    .cin(pp_0_11_5),
    .sum(pp_1_11_4),
    .cout(pp_1_12_1)
  );

  MG_FA fa_0_11_2(
    .a(pp_0_11_6),
    .b(pp_0_11_7),
    .cin(pp_0_11_8),
    .sum(pp_1_11_5),
    .cout(pp_1_12_2)
  );

  assign pp_1_11_6 = pp_0_11_9;
  assign pp_1_11_7 = pp_0_11_10;
  assign pp_1_11_8 = pp_0_11_11;
  MG_FA fa_0_12_0(
    .a(pp_0_12_0),
    .b(pp_0_12_1),
    .cin(pp_0_12_2),
    .sum(pp_1_12_3),
    .cout(pp_1_13_0)
  );

  MG_FA fa_0_12_1(
    .a(pp_0_12_3),
    .b(pp_0_12_4),
    .cin(pp_0_12_5),
    .sum(pp_1_12_4),
    .cout(pp_1_13_1)
  );

  MG_FA fa_0_12_2(
    .a(pp_0_12_6),
    .b(pp_0_12_7),
    .cin(pp_0_12_8),
    .sum(pp_1_12_5),
    .cout(pp_1_13_2)
  );

  MG_HA ha_0_12_3(
    .a(pp_0_12_9),
    .b(pp_0_12_10),
    .sum(pp_1_12_6),
    .cout(pp_1_13_3)
  );

  assign pp_1_12_7 = pp_0_12_11;
  assign pp_1_12_8 = pp_0_12_12;
  MG_FA fa_0_13_0(
    .a(pp_0_13_0),
    .b(pp_0_13_1),
    .cin(pp_0_13_2),
    .sum(pp_1_13_4),
    .cout(pp_1_14_0)
  );

  MG_FA fa_0_13_1(
    .a(pp_0_13_3),
    .b(pp_0_13_4),
    .cin(pp_0_13_5),
    .sum(pp_1_13_5),
    .cout(pp_1_14_1)
  );

  MG_FA fa_0_13_2(
    .a(pp_0_13_6),
    .b(pp_0_13_7),
    .cin(pp_0_13_8),
    .sum(pp_1_13_6),
    .cout(pp_1_14_2)
  );

  MG_FA fa_0_13_3(
    .a(pp_0_13_9),
    .b(pp_0_13_10),
    .cin(pp_0_13_11),
    .sum(pp_1_13_7),
    .cout(pp_1_14_3)
  );

  MG_HA ha_0_13_4(
    .a(pp_0_13_12),
    .b(pp_0_13_13),
    .sum(pp_1_13_8),
    .cout(pp_1_14_4)
  );

  assign pp_1_14_5 = pp_0_14_0;
  assign pp_1_14_6 = pp_0_14_1;
  assign pp_1_14_7 = pp_0_14_2;
  assign pp_1_14_8 = pp_0_14_3;
  assign pp_1_14_9 = pp_0_14_4;
  assign pp_1_14_10 = pp_0_14_5;
  assign pp_1_14_11 = pp_0_14_6;
  assign pp_1_14_12 = pp_0_14_7;
  assign pp_1_14_13 = pp_0_14_8;
  assign pp_1_14_14 = pp_0_14_9;
  assign pp_1_14_15 = pp_0_14_10;
  assign pp_1_14_16 = pp_0_14_11;
  assign pp_1_14_17 = pp_0_14_12;
  assign pp_1_14_18 = pp_0_14_13;
  assign pp_1_14_19 = pp_0_14_14;
  MG_FA fa_0_15_0(
    .a(pp_0_15_0),
    .b(pp_0_15_1),
    .cin(pp_0_15_2),
    .sum(pp_1_15_0),
    .cout(pp_1_16_0)
  );

  MG_FA fa_0_15_1(
    .a(pp_0_15_3),
    .b(pp_0_15_4),
    .cin(pp_0_15_5),
    .sum(pp_1_15_1),
    .cout(pp_1_16_1)
  );

  MG_FA fa_0_15_2(
    .a(pp_0_15_6),
    .b(pp_0_15_7),
    .cin(pp_0_15_8),
    .sum(pp_1_15_2),
    .cout(pp_1_16_2)
  );

  MG_FA fa_0_15_3(
    .a(pp_0_15_9),
    .b(pp_0_15_10),
    .cin(pp_0_15_11),
    .sum(pp_1_15_3),
    .cout(pp_1_16_3)
  );

  MG_FA fa_0_15_4(
    .a(pp_0_15_12),
    .b(pp_0_15_13),
    .cin(pp_0_15_14),
    .sum(pp_1_15_4),
    .cout(pp_1_16_4)
  );

  assign pp_1_15_5 = pp_0_15_15;
  assign pp_1_16_5 = pp_0_16_0;
  assign pp_1_16_6 = pp_0_16_1;
  assign pp_1_16_7 = pp_0_16_2;
  assign pp_1_16_8 = pp_0_16_3;
  assign pp_1_16_9 = pp_0_16_4;
  assign pp_1_16_10 = pp_0_16_5;
  assign pp_1_16_11 = pp_0_16_6;
  assign pp_1_16_12 = pp_0_16_7;
  assign pp_1_16_13 = pp_0_16_8;
  assign pp_1_16_14 = pp_0_16_9;
  assign pp_1_16_15 = pp_0_16_10;
  assign pp_1_16_16 = pp_0_16_11;
  assign pp_1_16_17 = pp_0_16_12;
  assign pp_1_16_18 = pp_0_16_13;
  assign pp_1_16_19 = pp_0_16_14;
  assign pp_1_16_20 = pp_0_16_15;
  MG_FA fa_0_17_0(
    .a(pp_0_17_0),
    .b(pp_0_17_1),
    .cin(pp_0_17_2),
    .sum(pp_1_17_0),
    .cout(pp_1_18_0)
  );

  MG_FA fa_0_17_1(
    .a(pp_0_17_3),
    .b(pp_0_17_4),
    .cin(pp_0_17_5),
    .sum(pp_1_17_1),
    .cout(pp_1_18_1)
  );

  MG_FA fa_0_17_2(
    .a(pp_0_17_6),
    .b(pp_0_17_7),
    .cin(pp_0_17_8),
    .sum(pp_1_17_2),
    .cout(pp_1_18_2)
  );

  MG_FA fa_0_17_3(
    .a(pp_0_17_9),
    .b(pp_0_17_10),
    .cin(pp_0_17_11),
    .sum(pp_1_17_3),
    .cout(pp_1_18_3)
  );

  assign pp_1_17_4 = pp_0_17_12;
  assign pp_1_17_5 = pp_0_17_13;
  MG_FA fa_0_18_0(
    .a(pp_0_18_0),
    .b(pp_0_18_1),
    .cin(pp_0_18_2),
    .sum(pp_1_18_4),
    .cout(pp_1_19_0)
  );

  MG_FA fa_0_18_1(
    .a(pp_0_18_3),
    .b(pp_0_18_4),
    .cin(pp_0_18_5),
    .sum(pp_1_18_5),
    .cout(pp_1_19_1)
  );

  MG_FA fa_0_18_2(
    .a(pp_0_18_6),
    .b(pp_0_18_7),
    .cin(pp_0_18_8),
    .sum(pp_1_18_6),
    .cout(pp_1_19_2)
  );

  MG_FA fa_0_18_3(
    .a(pp_0_18_9),
    .b(pp_0_18_10),
    .cin(pp_0_18_11),
    .sum(pp_1_18_7),
    .cout(pp_1_19_3)
  );

  assign pp_1_18_8 = pp_0_18_12;
  MG_FA fa_0_19_0(
    .a(pp_0_19_0),
    .b(pp_0_19_1),
    .cin(pp_0_19_2),
    .sum(pp_1_19_4),
    .cout(pp_1_20_0)
  );

  MG_FA fa_0_19_1(
    .a(pp_0_19_3),
    .b(pp_0_19_4),
    .cin(pp_0_19_5),
    .sum(pp_1_19_5),
    .cout(pp_1_20_1)
  );

  MG_FA fa_0_19_2(
    .a(pp_0_19_6),
    .b(pp_0_19_7),
    .cin(pp_0_19_8),
    .sum(pp_1_19_6),
    .cout(pp_1_20_2)
  );

  MG_FA fa_0_19_3(
    .a(pp_0_19_9),
    .b(pp_0_19_10),
    .cin(pp_0_19_11),
    .sum(pp_1_19_7),
    .cout(pp_1_20_3)
  );

  MG_FA fa_0_20_0(
    .a(pp_0_20_0),
    .b(pp_0_20_1),
    .cin(pp_0_20_2),
    .sum(pp_1_20_4),
    .cout(pp_1_21_0)
  );

  MG_FA fa_0_20_1(
    .a(pp_0_20_3),
    .b(pp_0_20_4),
    .cin(pp_0_20_5),
    .sum(pp_1_20_5),
    .cout(pp_1_21_1)
  );

  MG_FA fa_0_20_2(
    .a(pp_0_20_6),
    .b(pp_0_20_7),
    .cin(pp_0_20_8),
    .sum(pp_1_20_6),
    .cout(pp_1_21_2)
  );

  assign pp_1_20_7 = pp_0_20_9;
  assign pp_1_20_8 = pp_0_20_10;
  MG_FA fa_0_21_0(
    .a(pp_0_21_0),
    .b(pp_0_21_1),
    .cin(pp_0_21_2),
    .sum(pp_1_21_3),
    .cout(pp_1_22_0)
  );

  MG_FA fa_0_21_1(
    .a(pp_0_21_3),
    .b(pp_0_21_4),
    .cin(pp_0_21_5),
    .sum(pp_1_21_4),
    .cout(pp_1_22_1)
  );

  MG_FA fa_0_21_2(
    .a(pp_0_21_6),
    .b(pp_0_21_7),
    .cin(pp_0_21_8),
    .sum(pp_1_21_5),
    .cout(pp_1_22_2)
  );

  assign pp_1_21_6 = pp_0_21_9;
  MG_FA fa_0_22_0(
    .a(pp_0_22_0),
    .b(pp_0_22_1),
    .cin(pp_0_22_2),
    .sum(pp_1_22_3),
    .cout(pp_1_23_0)
  );

  MG_FA fa_0_22_1(
    .a(pp_0_22_3),
    .b(pp_0_22_4),
    .cin(pp_0_22_5),
    .sum(pp_1_22_4),
    .cout(pp_1_23_1)
  );

  MG_FA fa_0_22_2(
    .a(pp_0_22_6),
    .b(pp_0_22_7),
    .cin(pp_0_22_8),
    .sum(pp_1_22_5),
    .cout(pp_1_23_2)
  );

  assign pp_1_23_3 = pp_0_23_0;
  assign pp_1_23_4 = pp_0_23_1;
  assign pp_1_23_5 = pp_0_23_2;
  assign pp_1_23_6 = pp_0_23_3;
  assign pp_1_23_7 = pp_0_23_4;
  assign pp_1_23_8 = pp_0_23_5;
  assign pp_1_23_9 = pp_0_23_6;
  assign pp_1_23_10 = pp_0_23_7;
  MG_FA fa_0_24_0(
    .a(pp_0_24_0),
    .b(pp_0_24_1),
    .cin(pp_0_24_2),
    .sum(pp_1_24_0),
    .cout(pp_1_25_0)
  );

  assign pp_1_24_1 = pp_0_24_3;
  assign pp_1_24_2 = pp_0_24_4;
  assign pp_1_24_3 = pp_0_24_5;
  assign pp_1_24_4 = pp_0_24_6;
  MG_FA fa_0_25_0(
    .a(pp_0_25_0),
    .b(pp_0_25_1),
    .cin(pp_0_25_2),
    .sum(pp_1_25_1),
    .cout(pp_1_26_0)
  );

  MG_FA fa_0_25_1(
    .a(pp_0_25_3),
    .b(pp_0_25_4),
    .cin(pp_0_25_5),
    .sum(pp_1_25_2),
    .cout(pp_1_26_1)
  );

  assign pp_1_26_2 = pp_0_26_0;
  assign pp_1_26_3 = pp_0_26_1;
  assign pp_1_26_4 = pp_0_26_2;
  assign pp_1_26_5 = pp_0_26_3;
  assign pp_1_26_6 = pp_0_26_4;
  assign pp_1_27_0 = pp_0_27_0;
  assign pp_1_27_1 = pp_0_27_1;
  assign pp_1_27_2 = pp_0_27_2;
  assign pp_1_27_3 = pp_0_27_3;
  MG_FA fa_0_28_0(
    .a(pp_0_28_0),
    .b(pp_0_28_1),
    .cin(pp_0_28_2),
    .sum(pp_1_28_0),
    .cout(pp_1_29_0)
  );

  assign pp_1_29_1 = pp_0_29_0;
  assign pp_1_29_2 = pp_0_29_1;
  assign pp_1_30_0 = pp_0_30_0;
  assign pp_1_31_0 = pp_0_31_0;
  assign pp_2_0_0 = pp_1_0_0;
  assign pp_2_1_0 = pp_1_1_0;
  assign pp_2_1_1 = pp_1_1_1;
  assign pp_2_2_0 = pp_1_2_0;
  assign pp_2_2_1 = pp_1_2_1;
  assign pp_2_2_2 = pp_1_2_2;
  MG_FA fa_1_3_0(
    .a(pp_1_3_0),
    .b(pp_1_3_1),
    .cin(pp_1_3_2),
    .sum(pp_2_3_0),
    .cout(pp_2_4_0)
  );

  assign pp_2_3_1 = pp_1_3_3;
  MG_FA fa_1_4_0(
    .a(pp_1_4_0),
    .b(pp_1_4_1),
    .cin(pp_1_4_2),
    .sum(pp_2_4_1),
    .cout(pp_2_5_0)
  );

  MG_FA fa_1_5_0(
    .a(pp_1_5_0),
    .b(pp_1_5_1),
    .cin(pp_1_5_2),
    .sum(pp_2_5_1),
    .cout(pp_2_6_0)
  );

  MG_FA fa_1_6_0(
    .a(pp_1_6_0),
    .b(pp_1_6_1),
    .cin(pp_1_6_2),
    .sum(pp_2_6_1),
    .cout(pp_2_7_0)
  );

  MG_FA fa_1_6_1(
    .a(pp_1_6_3),
    .b(pp_1_6_4),
    .cin(pp_1_6_5),
    .sum(pp_2_6_2),
    .cout(pp_2_7_1)
  );

  MG_FA fa_1_6_2(
    .a(pp_1_6_6),
    .b(pp_1_6_7),
    .cin(pp_1_6_8),
    .sum(pp_2_6_3),
    .cout(pp_2_7_2)
  );

  MG_FA fa_1_7_0(
    .a(pp_1_7_0),
    .b(pp_1_7_1),
    .cin(pp_1_7_2),
    .sum(pp_2_7_3),
    .cout(pp_2_8_0)
  );

  MG_FA fa_1_8_0(
    .a(pp_1_8_0),
    .b(pp_1_8_1),
    .cin(pp_1_8_2),
    .sum(pp_2_8_1),
    .cout(pp_2_9_0)
  );

  MG_FA fa_1_8_1(
    .a(pp_1_8_3),
    .b(pp_1_8_4),
    .cin(pp_1_8_5),
    .sum(pp_2_8_2),
    .cout(pp_2_9_1)
  );

  MG_FA fa_1_8_2(
    .a(pp_1_8_6),
    .b(pp_1_8_7),
    .cin(pp_1_8_8),
    .sum(pp_2_8_3),
    .cout(pp_2_9_2)
  );

  MG_FA fa_1_8_3(
    .a(pp_1_8_9),
    .b(pp_1_8_10),
    .cin(pp_1_8_11),
    .sum(pp_2_8_4),
    .cout(pp_2_9_3)
  );

  MG_FA fa_1_9_0(
    .a(pp_1_9_0),
    .b(pp_1_9_1),
    .cin(pp_1_9_2),
    .sum(pp_2_9_4),
    .cout(pp_2_10_0)
  );

  MG_FA fa_1_9_1(
    .a(pp_1_9_3),
    .b(pp_1_9_4),
    .cin(pp_1_9_5),
    .sum(pp_2_9_5),
    .cout(pp_2_10_1)
  );

  MG_FA fa_1_9_2(
    .a(pp_1_9_6),
    .b(pp_1_9_7),
    .cin(pp_1_9_8),
    .sum(pp_2_9_6),
    .cout(pp_2_10_2)
  );

  assign pp_2_9_7 = pp_1_9_9;
  MG_FA fa_1_10_0(
    .a(pp_1_10_0),
    .b(pp_1_10_1),
    .cin(pp_1_10_2),
    .sum(pp_2_10_3),
    .cout(pp_2_11_0)
  );

  assign pp_2_10_4 = pp_1_10_3;
  assign pp_2_10_5 = pp_1_10_4;
  MG_FA fa_1_11_0(
    .a(pp_1_11_0),
    .b(pp_1_11_1),
    .cin(pp_1_11_2),
    .sum(pp_2_11_1),
    .cout(pp_2_12_0)
  );

  MG_FA fa_1_11_1(
    .a(pp_1_11_3),
    .b(pp_1_11_4),
    .cin(pp_1_11_5),
    .sum(pp_2_11_2),
    .cout(pp_2_12_1)
  );

  MG_FA fa_1_11_2(
    .a(pp_1_11_6),
    .b(pp_1_11_7),
    .cin(pp_1_11_8),
    .sum(pp_2_11_3),
    .cout(pp_2_12_2)
  );

  MG_FA fa_1_12_0(
    .a(pp_1_12_0),
    .b(pp_1_12_1),
    .cin(pp_1_12_2),
    .sum(pp_2_12_3),
    .cout(pp_2_13_0)
  );

  MG_FA fa_1_12_1(
    .a(pp_1_12_3),
    .b(pp_1_12_4),
    .cin(pp_1_12_5),
    .sum(pp_2_12_4),
    .cout(pp_2_13_1)
  );

  MG_FA fa_1_12_2(
    .a(pp_1_12_6),
    .b(pp_1_12_7),
    .cin(pp_1_12_8),
    .sum(pp_2_12_5),
    .cout(pp_2_13_2)
  );

  MG_FA fa_1_13_0(
    .a(pp_1_13_0),
    .b(pp_1_13_1),
    .cin(pp_1_13_2),
    .sum(pp_2_13_3),
    .cout(pp_2_14_0)
  );

  MG_FA fa_1_13_1(
    .a(pp_1_13_3),
    .b(pp_1_13_4),
    .cin(pp_1_13_5),
    .sum(pp_2_13_4),
    .cout(pp_2_14_1)
  );

  MG_FA fa_1_13_2(
    .a(pp_1_13_6),
    .b(pp_1_13_7),
    .cin(pp_1_13_8),
    .sum(pp_2_13_5),
    .cout(pp_2_14_2)
  );

  MG_FA fa_1_14_0(
    .a(pp_1_14_0),
    .b(pp_1_14_1),
    .cin(pp_1_14_2),
    .sum(pp_2_14_3),
    .cout(pp_2_15_0)
  );

  MG_FA fa_1_14_1(
    .a(pp_1_14_3),
    .b(pp_1_14_4),
    .cin(pp_1_14_5),
    .sum(pp_2_14_4),
    .cout(pp_2_15_1)
  );

  MG_FA fa_1_14_2(
    .a(pp_1_14_6),
    .b(pp_1_14_7),
    .cin(pp_1_14_8),
    .sum(pp_2_14_5),
    .cout(pp_2_15_2)
  );

  MG_FA fa_1_14_3(
    .a(pp_1_14_9),
    .b(pp_1_14_10),
    .cin(pp_1_14_11),
    .sum(pp_2_14_6),
    .cout(pp_2_15_3)
  );

  MG_FA fa_1_14_4(
    .a(pp_1_14_12),
    .b(pp_1_14_13),
    .cin(pp_1_14_14),
    .sum(pp_2_14_7),
    .cout(pp_2_15_4)
  );

  MG_FA fa_1_14_5(
    .a(pp_1_14_15),
    .b(pp_1_14_16),
    .cin(pp_1_14_17),
    .sum(pp_2_14_8),
    .cout(pp_2_15_5)
  );

  MG_HA ha_1_14_6(
    .a(pp_1_14_18),
    .b(pp_1_14_19),
    .sum(pp_2_14_9),
    .cout(pp_2_15_6)
  );

  MG_FA fa_1_15_0(
    .a(pp_1_15_0),
    .b(pp_1_15_1),
    .cin(pp_1_15_2),
    .sum(pp_2_15_7),
    .cout(pp_2_16_0)
  );

  MG_FA fa_1_15_1(
    .a(pp_1_15_3),
    .b(pp_1_15_4),
    .cin(pp_1_15_5),
    .sum(pp_2_15_8),
    .cout(pp_2_16_1)
  );

  MG_FA fa_1_16_0(
    .a(pp_1_16_0),
    .b(pp_1_16_1),
    .cin(pp_1_16_2),
    .sum(pp_2_16_2),
    .cout(pp_2_17_0)
  );

  MG_FA fa_1_16_1(
    .a(pp_1_16_3),
    .b(pp_1_16_4),
    .cin(pp_1_16_5),
    .sum(pp_2_16_3),
    .cout(pp_2_17_1)
  );

  MG_FA fa_1_16_2(
    .a(pp_1_16_6),
    .b(pp_1_16_7),
    .cin(pp_1_16_8),
    .sum(pp_2_16_4),
    .cout(pp_2_17_2)
  );

  MG_FA fa_1_16_3(
    .a(pp_1_16_9),
    .b(pp_1_16_10),
    .cin(pp_1_16_11),
    .sum(pp_2_16_5),
    .cout(pp_2_17_3)
  );

  MG_FA fa_1_16_4(
    .a(pp_1_16_12),
    .b(pp_1_16_13),
    .cin(pp_1_16_14),
    .sum(pp_2_16_6),
    .cout(pp_2_17_4)
  );

  MG_FA fa_1_16_5(
    .a(pp_1_16_15),
    .b(pp_1_16_16),
    .cin(pp_1_16_17),
    .sum(pp_2_16_7),
    .cout(pp_2_17_5)
  );

  MG_FA fa_1_16_6(
    .a(pp_1_16_18),
    .b(pp_1_16_19),
    .cin(pp_1_16_20),
    .sum(pp_2_16_8),
    .cout(pp_2_17_6)
  );

  MG_FA fa_1_17_0(
    .a(pp_1_17_0),
    .b(pp_1_17_1),
    .cin(pp_1_17_2),
    .sum(pp_2_17_7),
    .cout(pp_2_18_0)
  );

  MG_FA fa_1_17_1(
    .a(pp_1_17_3),
    .b(pp_1_17_4),
    .cin(pp_1_17_5),
    .sum(pp_2_17_8),
    .cout(pp_2_18_1)
  );

  MG_FA fa_1_18_0(
    .a(pp_1_18_0),
    .b(pp_1_18_1),
    .cin(pp_1_18_2),
    .sum(pp_2_18_2),
    .cout(pp_2_19_0)
  );

  MG_FA fa_1_18_1(
    .a(pp_1_18_3),
    .b(pp_1_18_4),
    .cin(pp_1_18_5),
    .sum(pp_2_18_3),
    .cout(pp_2_19_1)
  );

  MG_FA fa_1_18_2(
    .a(pp_1_18_6),
    .b(pp_1_18_7),
    .cin(pp_1_18_8),
    .sum(pp_2_18_4),
    .cout(pp_2_19_2)
  );

  MG_FA fa_1_19_0(
    .a(pp_1_19_0),
    .b(pp_1_19_1),
    .cin(pp_1_19_2),
    .sum(pp_2_19_3),
    .cout(pp_2_20_0)
  );

  MG_FA fa_1_19_1(
    .a(pp_1_19_3),
    .b(pp_1_19_4),
    .cin(pp_1_19_5),
    .sum(pp_2_19_4),
    .cout(pp_2_20_1)
  );

  assign pp_2_19_5 = pp_1_19_6;
  assign pp_2_19_6 = pp_1_19_7;
  MG_FA fa_1_20_0(
    .a(pp_1_20_0),
    .b(pp_1_20_1),
    .cin(pp_1_20_2),
    .sum(pp_2_20_2),
    .cout(pp_2_21_0)
  );

  MG_FA fa_1_20_1(
    .a(pp_1_20_3),
    .b(pp_1_20_4),
    .cin(pp_1_20_5),
    .sum(pp_2_20_3),
    .cout(pp_2_21_1)
  );

  MG_FA fa_1_20_2(
    .a(pp_1_20_6),
    .b(pp_1_20_7),
    .cin(pp_1_20_8),
    .sum(pp_2_20_4),
    .cout(pp_2_21_2)
  );

  MG_FA fa_1_21_0(
    .a(pp_1_21_0),
    .b(pp_1_21_1),
    .cin(pp_1_21_2),
    .sum(pp_2_21_3),
    .cout(pp_2_22_0)
  );

  MG_FA fa_1_21_1(
    .a(pp_1_21_3),
    .b(pp_1_21_4),
    .cin(pp_1_21_5),
    .sum(pp_2_21_4),
    .cout(pp_2_22_1)
  );

  assign pp_2_21_5 = pp_1_21_6;
  MG_FA fa_1_22_0(
    .a(pp_1_22_0),
    .b(pp_1_22_1),
    .cin(pp_1_22_2),
    .sum(pp_2_22_2),
    .cout(pp_2_23_0)
  );

  MG_FA fa_1_22_1(
    .a(pp_1_22_3),
    .b(pp_1_22_4),
    .cin(pp_1_22_5),
    .sum(pp_2_22_3),
    .cout(pp_2_23_1)
  );

  MG_FA fa_1_23_0(
    .a(pp_1_23_0),
    .b(pp_1_23_1),
    .cin(pp_1_23_2),
    .sum(pp_2_23_2),
    .cout(pp_2_24_0)
  );

  MG_FA fa_1_23_1(
    .a(pp_1_23_3),
    .b(pp_1_23_4),
    .cin(pp_1_23_5),
    .sum(pp_2_23_3),
    .cout(pp_2_24_1)
  );

  MG_FA fa_1_23_2(
    .a(pp_1_23_6),
    .b(pp_1_23_7),
    .cin(pp_1_23_8),
    .sum(pp_2_23_4),
    .cout(pp_2_24_2)
  );

  assign pp_2_23_5 = pp_1_23_9;
  assign pp_2_23_6 = pp_1_23_10;
  MG_FA fa_1_24_0(
    .a(pp_1_24_0),
    .b(pp_1_24_1),
    .cin(pp_1_24_2),
    .sum(pp_2_24_3),
    .cout(pp_2_25_0)
  );

  assign pp_2_24_4 = pp_1_24_3;
  assign pp_2_24_5 = pp_1_24_4;
  MG_FA fa_1_25_0(
    .a(pp_1_25_0),
    .b(pp_1_25_1),
    .cin(pp_1_25_2),
    .sum(pp_2_25_1),
    .cout(pp_2_26_0)
  );

  MG_FA fa_1_26_0(
    .a(pp_1_26_0),
    .b(pp_1_26_1),
    .cin(pp_1_26_2),
    .sum(pp_2_26_1),
    .cout(pp_2_27_0)
  );

  MG_FA fa_1_26_1(
    .a(pp_1_26_3),
    .b(pp_1_26_4),
    .cin(pp_1_26_5),
    .sum(pp_2_26_2),
    .cout(pp_2_27_1)
  );

  assign pp_2_26_3 = pp_1_26_6;
  MG_FA fa_1_27_0(
    .a(pp_1_27_0),
    .b(pp_1_27_1),
    .cin(pp_1_27_2),
    .sum(pp_2_27_2),
    .cout(pp_2_28_0)
  );

  assign pp_2_27_3 = pp_1_27_3;
  assign pp_2_28_1 = pp_1_28_0;
  MG_FA fa_1_29_0(
    .a(pp_1_29_0),
    .b(pp_1_29_1),
    .cin(pp_1_29_2),
    .sum(pp_2_29_0),
    .cout(pp_2_30_0)
  );

  assign pp_2_30_1 = pp_1_30_0;
  assign pp_2_31_0 = pp_1_31_0;
  assign pp_3_0_0 = pp_2_0_0;
  assign pp_3_1_0 = pp_2_1_0;
  assign pp_3_1_1 = pp_2_1_1;
  assign pp_3_2_0 = pp_2_2_0;
  assign pp_3_2_1 = pp_2_2_1;
  assign pp_3_2_2 = pp_2_2_2;
  assign pp_3_3_0 = pp_2_3_0;
  assign pp_3_3_1 = pp_2_3_1;
  assign pp_3_4_0 = pp_2_4_0;
  assign pp_3_4_1 = pp_2_4_1;
  assign pp_3_5_0 = pp_2_5_0;
  assign pp_3_5_1 = pp_2_5_1;
  assign pp_3_6_0 = pp_2_6_0;
  assign pp_3_6_1 = pp_2_6_1;
  assign pp_3_6_2 = pp_2_6_2;
  assign pp_3_6_3 = pp_2_6_3;
  MG_FA fa_2_7_0(
    .a(pp_2_7_0),
    .b(pp_2_7_1),
    .cin(pp_2_7_2),
    .sum(pp_3_7_0),
    .cout(pp_3_8_0)
  );

  assign pp_3_7_1 = pp_2_7_3;
  assign pp_3_8_1 = pp_2_8_0;
  assign pp_3_8_2 = pp_2_8_1;
  assign pp_3_8_3 = pp_2_8_2;
  assign pp_3_8_4 = pp_2_8_3;
  assign pp_3_8_5 = pp_2_8_4;
  MG_FA fa_2_9_0(
    .a(pp_2_9_0),
    .b(pp_2_9_1),
    .cin(pp_2_9_2),
    .sum(pp_3_9_0),
    .cout(pp_3_10_0)
  );

  MG_FA fa_2_9_1(
    .a(pp_2_9_3),
    .b(pp_2_9_4),
    .cin(pp_2_9_5),
    .sum(pp_3_9_1),
    .cout(pp_3_10_1)
  );

  MG_HA ha_2_9_2(
    .a(pp_2_9_6),
    .b(pp_2_9_7),
    .sum(pp_3_9_2),
    .cout(pp_3_10_2)
  );

  MG_FA fa_2_10_0(
    .a(pp_2_10_0),
    .b(pp_2_10_1),
    .cin(pp_2_10_2),
    .sum(pp_3_10_3),
    .cout(pp_3_11_0)
  );

  MG_FA fa_2_10_1(
    .a(pp_2_10_3),
    .b(pp_2_10_4),
    .cin(pp_2_10_5),
    .sum(pp_3_10_4),
    .cout(pp_3_11_1)
  );

  MG_FA fa_2_11_0(
    .a(pp_2_11_0),
    .b(pp_2_11_1),
    .cin(pp_2_11_2),
    .sum(pp_3_11_2),
    .cout(pp_3_12_0)
  );

  assign pp_3_11_3 = pp_2_11_3;
  MG_FA fa_2_12_0(
    .a(pp_2_12_0),
    .b(pp_2_12_1),
    .cin(pp_2_12_2),
    .sum(pp_3_12_1),
    .cout(pp_3_13_0)
  );

  MG_FA fa_2_12_1(
    .a(pp_2_12_3),
    .b(pp_2_12_4),
    .cin(pp_2_12_5),
    .sum(pp_3_12_2),
    .cout(pp_3_13_1)
  );

  MG_FA fa_2_13_0(
    .a(pp_2_13_0),
    .b(pp_2_13_1),
    .cin(pp_2_13_2),
    .sum(pp_3_13_2),
    .cout(pp_3_14_0)
  );

  MG_FA fa_2_13_1(
    .a(pp_2_13_3),
    .b(pp_2_13_4),
    .cin(pp_2_13_5),
    .sum(pp_3_13_3),
    .cout(pp_3_14_1)
  );

  MG_FA fa_2_14_0(
    .a(pp_2_14_0),
    .b(pp_2_14_1),
    .cin(pp_2_14_2),
    .sum(pp_3_14_2),
    .cout(pp_3_15_0)
  );

  MG_FA fa_2_14_1(
    .a(pp_2_14_3),
    .b(pp_2_14_4),
    .cin(pp_2_14_5),
    .sum(pp_3_14_3),
    .cout(pp_3_15_1)
  );

  MG_FA fa_2_14_2(
    .a(pp_2_14_6),
    .b(pp_2_14_7),
    .cin(pp_2_14_8),
    .sum(pp_3_14_4),
    .cout(pp_3_15_2)
  );

  assign pp_3_14_5 = pp_2_14_9;
  MG_FA fa_2_15_0(
    .a(pp_2_15_0),
    .b(pp_2_15_1),
    .cin(pp_2_15_2),
    .sum(pp_3_15_3),
    .cout(pp_3_16_0)
  );

  MG_FA fa_2_15_1(
    .a(pp_2_15_3),
    .b(pp_2_15_4),
    .cin(pp_2_15_5),
    .sum(pp_3_15_4),
    .cout(pp_3_16_1)
  );

  MG_FA fa_2_15_2(
    .a(pp_2_15_6),
    .b(pp_2_15_7),
    .cin(pp_2_15_8),
    .sum(pp_3_15_5),
    .cout(pp_3_16_2)
  );

  MG_FA fa_2_16_0(
    .a(pp_2_16_0),
    .b(pp_2_16_1),
    .cin(pp_2_16_2),
    .sum(pp_3_16_3),
    .cout(pp_3_17_0)
  );

  MG_FA fa_2_16_1(
    .a(pp_2_16_3),
    .b(pp_2_16_4),
    .cin(pp_2_16_5),
    .sum(pp_3_16_4),
    .cout(pp_3_17_1)
  );

  MG_FA fa_2_16_2(
    .a(pp_2_16_6),
    .b(pp_2_16_7),
    .cin(pp_2_16_8),
    .sum(pp_3_16_5),
    .cout(pp_3_17_2)
  );

  MG_FA fa_2_17_0(
    .a(pp_2_17_0),
    .b(pp_2_17_1),
    .cin(pp_2_17_7),
    .sum(pp_3_17_3),
    .cout(pp_3_18_0)
  );

  MG_FA fa_2_17_1(
    .a(pp_2_17_3),
    .b(pp_2_17_4),
    .cin(pp_2_17_5),
    .sum(pp_3_17_4),
    .cout(pp_3_18_1)
  );

  MG_FA fa_2_17_2(
    .a(pp_2_17_6),
    .b(pp_2_17_2),
    .cin(pp_2_17_8),
    .sum(pp_3_17_5),
    .cout(pp_3_18_2)
  );

  MG_FA fa_2_18_0(
    .a(pp_2_18_0),
    .b(pp_2_18_1),
    .cin(pp_2_18_2),
    .sum(pp_3_18_3),
    .cout(pp_3_19_0)
  );

  assign pp_3_18_4 = pp_2_18_3;
  assign pp_3_18_5 = pp_2_18_4;
  MG_FA fa_2_19_0(
    .a(pp_2_19_0),
    .b(pp_2_19_1),
    .cin(pp_2_19_2),
    .sum(pp_3_19_1),
    .cout(pp_3_20_0)
  );

  assign pp_3_19_2 = pp_2_19_3;
  assign pp_3_19_3 = pp_2_19_4;
  assign pp_3_19_4 = pp_2_19_5;
  assign pp_3_19_5 = pp_2_19_6;
  MG_FA fa_2_20_0(
    .a(pp_2_20_0),
    .b(pp_2_20_1),
    .cin(pp_2_20_2),
    .sum(pp_3_20_1),
    .cout(pp_3_21_0)
  );

  assign pp_3_20_2 = pp_2_20_3;
  assign pp_3_20_3 = pp_2_20_4;
  MG_FA fa_2_21_0(
    .a(pp_2_21_0),
    .b(pp_2_21_1),
    .cin(pp_2_21_2),
    .sum(pp_3_21_1),
    .cout(pp_3_22_0)
  );

  MG_FA fa_2_21_1(
    .a(pp_2_21_3),
    .b(pp_2_21_4),
    .cin(pp_2_21_5),
    .sum(pp_3_21_2),
    .cout(pp_3_22_1)
  );

  assign pp_3_22_2 = pp_2_22_0;
  assign pp_3_22_3 = pp_2_22_1;
  assign pp_3_22_4 = pp_2_22_2;
  assign pp_3_22_5 = pp_2_22_3;
  MG_FA fa_2_23_0(
    .a(pp_2_23_0),
    .b(pp_2_23_1),
    .cin(pp_2_23_2),
    .sum(pp_3_23_0),
    .cout(pp_3_24_0)
  );

  MG_FA fa_2_23_1(
    .a(pp_2_23_3),
    .b(pp_2_23_4),
    .cin(pp_2_23_5),
    .sum(pp_3_23_1),
    .cout(pp_3_24_1)
  );

  assign pp_3_23_2 = pp_2_23_6;
  MG_FA fa_2_24_0(
    .a(pp_2_24_0),
    .b(pp_2_24_1),
    .cin(pp_2_24_2),
    .sum(pp_3_24_2),
    .cout(pp_3_25_0)
  );

  assign pp_3_24_3 = pp_2_24_3;
  assign pp_3_24_4 = pp_2_24_4;
  assign pp_3_24_5 = pp_2_24_5;
  assign pp_3_25_1 = pp_2_25_0;
  assign pp_3_25_2 = pp_2_25_1;
  assign pp_3_26_0 = pp_2_26_0;
  assign pp_3_26_1 = pp_2_26_1;
  assign pp_3_26_2 = pp_2_26_2;
  assign pp_3_26_3 = pp_2_26_3;
  MG_FA fa_2_27_0(
    .a(pp_2_27_0),
    .b(pp_2_27_1),
    .cin(pp_2_27_2),
    .sum(pp_3_27_0),
    .cout(pp_3_28_0)
  );

  assign pp_3_27_1 = pp_2_27_3;
  assign pp_3_28_1 = pp_2_28_0;
  assign pp_3_28_2 = pp_2_28_1;
  assign pp_3_29_0 = pp_2_29_0;
  assign pp_3_30_0 = pp_2_30_0;
  assign pp_3_30_1 = pp_2_30_1;
  assign pp_3_31_0 = pp_2_31_0;
  assign pp_4_0_0 = pp_3_0_0;
  assign pp_4_1_0 = pp_3_1_0;
  assign pp_4_1_1 = pp_3_1_1;
  assign pp_4_2_0 = pp_3_2_0;
  assign pp_4_2_1 = pp_3_2_1;
  assign pp_4_2_2 = pp_3_2_2;
  assign pp_4_3_0 = pp_3_3_0;
  assign pp_4_3_1 = pp_3_3_1;
  assign pp_4_4_0 = pp_3_4_0;
  assign pp_4_4_1 = pp_3_4_1;
  assign pp_4_5_0 = pp_3_5_0;
  assign pp_4_5_1 = pp_3_5_1;
  MG_FA fa_3_6_0(
    .a(pp_3_6_0),
    .b(pp_3_6_1),
    .cin(pp_3_6_2),
    .sum(pp_4_6_0),
    .cout(pp_4_7_0)
  );

  assign pp_4_6_1 = pp_3_6_3;
  assign pp_4_7_1 = pp_3_7_0;
  assign pp_4_7_2 = pp_3_7_1;
  MG_FA fa_3_8_0(
    .a(pp_3_8_0),
    .b(pp_3_8_1),
    .cin(pp_3_8_2),
    .sum(pp_4_8_0),
    .cout(pp_4_9_0)
  );

  MG_FA fa_3_8_1(
    .a(pp_3_8_3),
    .b(pp_3_8_4),
    .cin(pp_3_8_5),
    .sum(pp_4_8_1),
    .cout(pp_4_9_1)
  );

  MG_FA fa_3_9_0(
    .a(pp_3_9_0),
    .b(pp_3_9_1),
    .cin(pp_3_9_2),
    .sum(pp_4_9_2),
    .cout(pp_4_10_0)
  );

  MG_FA fa_3_10_0(
    .a(pp_3_10_0),
    .b(pp_3_10_1),
    .cin(pp_3_10_2),
    .sum(pp_4_10_1),
    .cout(pp_4_11_0)
  );

  MG_HA ha_3_10_1(
    .a(pp_3_10_3),
    .b(pp_3_10_4),
    .sum(pp_4_10_2),
    .cout(pp_4_11_1)
  );

  assign pp_4_11_2 = pp_3_11_0;
  assign pp_4_11_3 = pp_3_11_1;
  assign pp_4_11_4 = pp_3_11_2;
  assign pp_4_11_5 = pp_3_11_3;
  assign pp_4_12_0 = pp_3_12_0;
  assign pp_4_12_1 = pp_3_12_1;
  assign pp_4_12_2 = pp_3_12_2;
  assign pp_4_13_0 = pp_3_13_0;
  assign pp_4_13_1 = pp_3_13_1;
  assign pp_4_13_2 = pp_3_13_2;
  assign pp_4_13_3 = pp_3_13_3;
  MG_FA fa_3_14_0(
    .a(pp_3_14_0),
    .b(pp_3_14_1),
    .cin(pp_3_14_2),
    .sum(pp_4_14_0),
    .cout(pp_4_15_0)
  );

  MG_FA fa_3_14_1(
    .a(pp_3_14_3),
    .b(pp_3_14_4),
    .cin(pp_3_14_5),
    .sum(pp_4_14_1),
    .cout(pp_4_15_1)
  );

  MG_FA fa_3_15_0(
    .a(pp_3_15_0),
    .b(pp_3_15_1),
    .cin(pp_3_15_2),
    .sum(pp_4_15_2),
    .cout(pp_4_16_0)
  );

  assign pp_4_15_3 = pp_3_15_3;
  assign pp_4_15_4 = pp_3_15_4;
  assign pp_4_15_5 = pp_3_15_5;
  MG_FA fa_3_16_0(
    .a(pp_3_16_0),
    .b(pp_3_16_1),
    .cin(pp_3_16_2),
    .sum(pp_4_16_1),
    .cout(pp_4_17_0)
  );

  MG_FA fa_3_16_1(
    .a(pp_3_16_3),
    .b(pp_3_16_4),
    .cin(pp_3_16_5),
    .sum(pp_4_16_2),
    .cout(pp_4_17_1)
  );

  MG_FA fa_3_17_0(
    .a(pp_3_17_0),
    .b(pp_3_17_1),
    .cin(pp_3_17_2),
    .sum(pp_4_17_2),
    .cout(pp_4_18_0)
  );

  MG_FA fa_3_17_1(
    .a(pp_3_17_3),
    .b(pp_3_17_4),
    .cin(pp_3_17_5),
    .sum(pp_4_17_3),
    .cout(pp_4_18_1)
  );

  MG_FA fa_3_18_0(
    .a(pp_3_18_0),
    .b(pp_3_18_1),
    .cin(pp_3_18_2),
    .sum(pp_4_18_2),
    .cout(pp_4_19_0)
  );

  MG_FA fa_3_18_1(
    .a(pp_3_18_3),
    .b(pp_3_18_4),
    .cin(pp_3_18_5),
    .sum(pp_4_18_3),
    .cout(pp_4_19_1)
  );

  MG_FA fa_3_19_0(
    .a(pp_3_19_0),
    .b(pp_3_19_1),
    .cin(pp_3_19_2),
    .sum(pp_4_19_2),
    .cout(pp_4_20_0)
  );

  MG_FA fa_3_19_1(
    .a(pp_3_19_3),
    .b(pp_3_19_4),
    .cin(pp_3_19_5),
    .sum(pp_4_19_3),
    .cout(pp_4_20_1)
  );

  assign pp_4_20_2 = pp_3_20_0;
  assign pp_4_20_3 = pp_3_20_1;
  assign pp_4_20_4 = pp_3_20_2;
  assign pp_4_20_5 = pp_3_20_3;
  MG_FA fa_3_21_0(
    .a(pp_3_21_0),
    .b(pp_3_21_1),
    .cin(pp_3_21_2),
    .sum(pp_4_21_0),
    .cout(pp_4_22_0)
  );

  MG_FA fa_3_22_0(
    .a(pp_3_22_0),
    .b(pp_3_22_1),
    .cin(pp_3_22_2),
    .sum(pp_4_22_1),
    .cout(pp_4_23_0)
  );

  MG_FA fa_3_22_1(
    .a(pp_3_22_3),
    .b(pp_3_22_4),
    .cin(pp_3_22_5),
    .sum(pp_4_22_2),
    .cout(pp_4_23_1)
  );

  assign pp_4_23_2 = pp_3_23_0;
  assign pp_4_23_3 = pp_3_23_1;
  assign pp_4_23_4 = pp_3_23_2;
  MG_FA fa_3_24_0(
    .a(pp_3_24_0),
    .b(pp_3_24_1),
    .cin(pp_3_24_2),
    .sum(pp_4_24_0),
    .cout(pp_4_25_0)
  );

  MG_FA fa_3_24_1(
    .a(pp_3_24_3),
    .b(pp_3_24_4),
    .cin(pp_3_24_5),
    .sum(pp_4_24_1),
    .cout(pp_4_25_1)
  );

  MG_FA fa_3_25_0(
    .a(pp_3_25_0),
    .b(pp_3_25_1),
    .cin(pp_3_25_2),
    .sum(pp_4_25_2),
    .cout(pp_4_26_0)
  );

  MG_FA fa_3_26_0(
    .a(pp_3_26_0),
    .b(pp_3_26_1),
    .cin(pp_3_26_2),
    .sum(pp_4_26_1),
    .cout(pp_4_27_0)
  );

  assign pp_4_26_2 = pp_3_26_3;
  assign pp_4_27_1 = pp_3_27_0;
  assign pp_4_27_2 = pp_3_27_1;
  assign pp_4_28_0 = pp_3_28_0;
  assign pp_4_28_1 = pp_3_28_1;
  assign pp_4_28_2 = pp_3_28_2;
  assign pp_4_29_0 = pp_3_29_0;
  assign pp_4_30_0 = pp_3_30_0;
  assign pp_4_30_1 = pp_3_30_1;
  assign pp_4_31_0 = pp_3_31_0;
  assign pp_5_0_0 = pp_4_0_0;
  assign pp_5_1_0 = pp_4_1_0;
  assign pp_5_1_1 = pp_4_1_1;
  assign pp_5_2_0 = pp_4_2_0;
  assign pp_5_2_1 = pp_4_2_1;
  assign pp_5_2_2 = pp_4_2_2;
  MG_HA ha_4_3_0(
    .a(pp_4_3_0),
    .b(pp_4_3_1),
    .sum(pp_5_3_0),
    .cout(pp_5_4_0)
  );

  MG_HA ha_4_4_0(
    .a(pp_4_4_0),
    .b(pp_4_4_1),
    .sum(pp_5_4_1),
    .cout(pp_5_5_0)
  );

  MG_HA ha_4_5_0(
    .a(pp_4_5_0),
    .b(pp_4_5_1),
    .sum(pp_5_5_1),
    .cout(pp_5_6_0)
  );

  MG_HA ha_4_6_0(
    .a(pp_4_6_0),
    .b(pp_4_6_1),
    .sum(pp_5_6_1),
    .cout(pp_5_7_0)
  );

  MG_FA fa_4_7_0(
    .a(pp_4_7_0),
    .b(pp_4_7_1),
    .cin(pp_4_7_2),
    .sum(pp_5_7_1),
    .cout(pp_5_8_0)
  );

  assign pp_5_8_1 = pp_4_8_0;
  assign pp_5_8_2 = pp_4_8_1;
  assign pp_5_9_0 = pp_4_9_0;
  assign pp_5_9_1 = pp_4_9_1;
  assign pp_5_9_2 = pp_4_9_2;
  MG_FA fa_4_10_0(
    .a(pp_4_10_0),
    .b(pp_4_10_1),
    .cin(pp_4_10_2),
    .sum(pp_5_10_0),
    .cout(pp_5_11_0)
  );

  MG_FA fa_4_11_0(
    .a(pp_4_11_0),
    .b(pp_4_11_1),
    .cin(pp_4_11_2),
    .sum(pp_5_11_1),
    .cout(pp_5_12_0)
  );

  MG_FA fa_4_11_1(
    .a(pp_4_11_3),
    .b(pp_4_11_4),
    .cin(pp_4_11_5),
    .sum(pp_5_11_2),
    .cout(pp_5_12_1)
  );

  MG_FA fa_4_12_0(
    .a(pp_4_12_0),
    .b(pp_4_12_1),
    .cin(pp_4_12_2),
    .sum(pp_5_12_2),
    .cout(pp_5_13_0)
  );

  MG_FA fa_4_13_0(
    .a(pp_4_13_0),
    .b(pp_4_13_1),
    .cin(pp_4_13_2),
    .sum(pp_5_13_1),
    .cout(pp_5_14_0)
  );

  assign pp_5_13_2 = pp_4_13_3;
  assign pp_5_14_1 = pp_4_14_0;
  assign pp_5_14_2 = pp_4_14_1;
  MG_FA fa_4_15_0(
    .a(pp_4_15_0),
    .b(pp_4_15_1),
    .cin(pp_4_15_2),
    .sum(pp_5_15_0),
    .cout(pp_5_16_0)
  );

  MG_FA fa_4_15_1(
    .a(pp_4_15_3),
    .b(pp_4_15_4),
    .cin(pp_4_15_5),
    .sum(pp_5_15_1),
    .cout(pp_5_16_1)
  );

  MG_FA fa_4_16_0(
    .a(pp_4_16_0),
    .b(pp_4_16_1),
    .cin(pp_4_16_2),
    .sum(pp_5_16_2),
    .cout(pp_5_17_0)
  );

  MG_FA fa_4_17_0(
    .a(pp_4_17_0),
    .b(pp_4_17_1),
    .cin(pp_4_17_2),
    .sum(pp_5_17_1),
    .cout(pp_5_18_0)
  );

  assign pp_5_17_2 = pp_4_17_3;
  MG_FA fa_4_18_0(
    .a(pp_4_18_0),
    .b(pp_4_18_1),
    .cin(pp_4_18_2),
    .sum(pp_5_18_1),
    .cout(pp_5_19_0)
  );

  assign pp_5_18_2 = pp_4_18_3;
  MG_FA fa_4_19_0(
    .a(pp_4_19_0),
    .b(pp_4_19_1),
    .cin(pp_4_19_2),
    .sum(pp_5_19_1),
    .cout(pp_5_20_0)
  );

  assign pp_5_19_2 = pp_4_19_3;
  MG_FA fa_4_20_0(
    .a(pp_4_20_0),
    .b(pp_4_20_1),
    .cin(pp_4_20_2),
    .sum(pp_5_20_1),
    .cout(pp_5_21_0)
  );

  MG_FA fa_4_20_1(
    .a(pp_4_20_3),
    .b(pp_4_20_4),
    .cin(pp_4_20_5),
    .sum(pp_5_20_2),
    .cout(pp_5_21_1)
  );

  assign pp_5_21_2 = pp_4_21_0;
  assign pp_5_22_0 = pp_4_22_0;
  assign pp_5_22_1 = pp_4_22_1;
  assign pp_5_22_2 = pp_4_22_2;
  MG_FA fa_4_23_0(
    .a(pp_4_23_0),
    .b(pp_4_23_1),
    .cin(pp_4_23_2),
    .sum(pp_5_23_0),
    .cout(pp_5_24_0)
  );

  assign pp_5_23_1 = pp_4_23_3;
  assign pp_5_23_2 = pp_4_23_4;
  assign pp_5_24_1 = pp_4_24_0;
  assign pp_5_24_2 = pp_4_24_1;
  MG_FA fa_4_25_0(
    .a(pp_4_25_0),
    .b(pp_4_25_1),
    .cin(pp_4_25_2),
    .sum(pp_5_25_0),
    .cout(pp_5_26_0)
  );

  assign pp_5_26_1 = pp_4_26_0;
  assign pp_5_26_2 = pp_4_26_1;
  assign pp_5_26_3 = pp_4_26_2;
  MG_FA fa_4_27_0(
    .a(pp_4_27_0),
    .b(pp_4_27_1),
    .cin(pp_4_27_2),
    .sum(pp_5_27_0),
    .cout(pp_5_28_0)
  );

  assign pp_5_28_1 = pp_4_28_0;
  assign pp_5_28_2 = pp_4_28_1;
  assign pp_5_28_3 = pp_4_28_2;
  assign pp_5_29_0 = pp_4_29_0;
  assign pp_5_30_0 = pp_4_30_0;
  assign pp_5_30_1 = pp_4_30_1;
  assign pp_5_31_0 = pp_4_31_0;
  assign pp_6_0_0 = pp_5_0_0;
  assign pp_6_1_0 = pp_5_1_0;
  assign pp_6_1_1 = pp_5_1_1;
  MG_HA ha_5_2_0(
    .a(pp_5_2_0),
    .b(pp_5_2_1),
    .sum(pp_6_2_0),
    .cout(pp_6_3_0)
  );

  assign pp_6_2_1 = pp_5_2_2;
  assign pp_6_3_1 = pp_5_3_0;
  assign pp_6_4_0 = pp_5_4_0;
  assign pp_6_4_1 = pp_5_4_1;
  assign pp_6_5_0 = pp_5_5_0;
  assign pp_6_5_1 = pp_5_5_1;
  assign pp_6_6_0 = pp_5_6_0;
  assign pp_6_6_1 = pp_5_6_1;
  assign pp_6_7_0 = pp_5_7_0;
  assign pp_6_7_1 = pp_5_7_1;
  MG_HA ha_5_8_0(
    .a(pp_5_8_0),
    .b(pp_5_8_1),
    .sum(pp_6_8_0),
    .cout(pp_6_9_0)
  );

  assign pp_6_8_1 = pp_5_8_2;
  MG_FA fa_5_9_0(
    .a(pp_5_9_0),
    .b(pp_5_9_1),
    .cin(pp_5_9_2),
    .sum(pp_6_9_1),
    .cout(pp_6_10_0)
  );

  assign pp_6_10_1 = pp_5_10_0;
  MG_HA ha_5_11_0(
    .a(pp_5_11_0),
    .b(pp_5_11_1),
    .sum(pp_6_11_0),
    .cout(pp_6_12_0)
  );

  assign pp_6_11_1 = pp_5_11_2;
  MG_FA fa_5_12_0(
    .a(pp_5_12_0),
    .b(pp_5_12_1),
    .cin(pp_5_12_2),
    .sum(pp_6_12_1),
    .cout(pp_6_13_0)
  );

  MG_FA fa_5_13_0(
    .a(pp_5_13_0),
    .b(pp_5_13_1),
    .cin(pp_5_13_2),
    .sum(pp_6_13_1),
    .cout(pp_6_14_0)
  );

  MG_FA fa_5_14_0(
    .a(pp_5_14_0),
    .b(pp_5_14_1),
    .cin(pp_5_14_2),
    .sum(pp_6_14_1),
    .cout(pp_6_15_0)
  );

  MG_HA ha_5_15_0(
    .a(pp_5_15_0),
    .b(pp_5_15_1),
    .sum(pp_6_15_1),
    .cout(pp_6_16_0)
  );

  MG_FA fa_5_16_0(
    .a(pp_5_16_0),
    .b(pp_5_16_1),
    .cin(pp_5_16_2),
    .sum(pp_6_16_1),
    .cout(pp_6_17_0)
  );

  MG_FA fa_5_17_0(
    .a(pp_5_17_0),
    .b(pp_5_17_1),
    .cin(pp_5_17_2),
    .sum(pp_6_17_1),
    .cout(pp_6_18_0)
  );

  MG_FA fa_5_18_0(
    .a(pp_5_18_0),
    .b(pp_5_18_1),
    .cin(pp_5_18_2),
    .sum(pp_6_18_1),
    .cout(pp_6_19_0)
  );

  MG_FA fa_5_19_0(
    .a(pp_5_19_0),
    .b(pp_5_19_1),
    .cin(pp_5_19_2),
    .sum(pp_6_19_1),
    .cout(pp_6_20_0)
  );

  MG_FA fa_5_20_0(
    .a(pp_5_20_0),
    .b(pp_5_20_1),
    .cin(pp_5_20_2),
    .sum(pp_6_20_1),
    .cout(pp_6_21_0)
  );

  MG_FA fa_5_21_0(
    .a(pp_5_21_0),
    .b(pp_5_21_1),
    .cin(pp_5_21_2),
    .sum(pp_6_21_1),
    .cout(pp_6_22_0)
  );

  MG_FA fa_5_22_0(
    .a(pp_5_22_0),
    .b(pp_5_22_1),
    .cin(pp_5_22_2),
    .sum(pp_6_22_1),
    .cout(pp_6_23_0)
  );

  MG_FA fa_5_23_0(
    .a(pp_5_23_0),
    .b(pp_5_23_1),
    .cin(pp_5_23_2),
    .sum(pp_6_23_1),
    .cout(pp_6_24_0)
  );

  MG_FA fa_5_24_0(
    .a(pp_5_24_0),
    .b(pp_5_24_1),
    .cin(pp_5_24_2),
    .sum(pp_6_24_1),
    .cout(pp_6_25_0)
  );

  assign pp_6_25_1 = pp_5_25_0;
  MG_FA fa_5_26_0(
    .a(pp_5_26_0),
    .b(pp_5_26_1),
    .cin(pp_5_26_2),
    .sum(pp_6_26_0),
    .cout(pp_6_27_0)
  );

  assign pp_6_26_1 = pp_5_26_3;
  assign pp_6_27_1 = pp_5_27_0;
  MG_FA fa_5_28_0(
    .a(pp_5_28_0),
    .b(pp_5_28_1),
    .cin(pp_5_28_2),
    .sum(pp_6_28_0),
    .cout(pp_6_29_0)
  );

  assign pp_6_28_1 = pp_5_28_3;
  assign pp_6_29_1 = pp_5_29_0;
  assign pp_6_30_0 = pp_5_30_0;
  assign pp_6_30_1 = pp_5_30_1;
  assign pp_6_31_0 = pp_5_31_0;
  wire [30:0] cta;
  wire [30:0] ctb;
  wire [30:0] cts;
  wire ctc;

  MG_CPA cpa(
 .a(cta), .b(ctb), .sum(cts), .cout(ctc)
  );

  assign cta[0] = pp_6_1_0;
  assign ctb[0] = pp_6_1_1;
  assign cta[1] = pp_6_2_0;
  assign ctb[1] = pp_6_2_1;
  assign cta[2] = pp_6_3_0;
  assign ctb[2] = pp_6_3_1;
  assign cta[3] = pp_6_4_0;
  assign ctb[3] = pp_6_4_1;
  assign cta[4] = pp_6_5_0;
  assign ctb[4] = pp_6_5_1;
  assign cta[5] = pp_6_6_0;
  assign ctb[5] = pp_6_6_1;
  assign cta[6] = pp_6_7_0;
  assign ctb[6] = pp_6_7_1;
  assign cta[7] = pp_6_8_0;
  assign ctb[7] = pp_6_8_1;
  assign cta[8] = pp_6_9_0;
  assign ctb[8] = pp_6_9_1;
  assign cta[9] = pp_6_10_0;
  assign ctb[9] = pp_6_10_1;
  assign cta[10] = pp_6_11_0;
  assign ctb[10] = pp_6_11_1;
  assign cta[11] = pp_6_12_0;
  assign ctb[11] = pp_6_12_1;
  assign cta[12] = pp_6_13_0;
  assign ctb[12] = pp_6_13_1;
  assign cta[13] = pp_6_14_0;
  assign ctb[13] = pp_6_14_1;
  assign cta[14] = pp_6_15_0;
  assign ctb[14] = pp_6_15_1;
  assign cta[15] = pp_6_16_0;
  assign ctb[15] = pp_6_16_1;
  assign cta[16] = pp_6_17_0;
  assign ctb[16] = pp_6_17_1;
  assign cta[17] = pp_6_18_0;
  assign ctb[17] = pp_6_18_1;
  assign cta[18] = pp_6_19_0;
  assign ctb[18] = pp_6_19_1;
  assign cta[19] = pp_6_20_0;
  assign ctb[19] = pp_6_20_1;
  assign cta[20] = pp_6_21_0;
  assign ctb[20] = pp_6_21_1;
  assign cta[21] = pp_6_22_0;
  assign ctb[21] = pp_6_22_1;
  assign cta[22] = pp_6_23_0;
  assign ctb[22] = pp_6_23_1;
  assign cta[23] = pp_6_24_0;
  assign ctb[23] = pp_6_24_1;
  assign cta[24] = pp_6_25_0;
  assign ctb[24] = pp_6_25_1;
  assign cta[25] = pp_6_26_0;
  assign ctb[25] = pp_6_26_1;
  assign cta[26] = pp_6_27_0;
  assign ctb[26] = pp_6_27_1;
  assign cta[27] = pp_6_28_0;
  assign ctb[27] = pp_6_28_1;
  assign cta[28] = pp_6_29_0;
  assign ctb[28] = pp_6_29_1;
  assign cta[29] = pp_6_30_0;
  assign ctb[29] = pp_6_30_1;
  assign cta[30] = pp_6_31_0;
  assign ctb[30] = 1'b0;
  assign product[0] = pp_6_0_0;
  assign product[31:1] = cts;
endmodule
