module MG_FA(
  input a,
  input b,
  input cin,
  output sum,
  output cout
);

  assign sum = (a ^ b) ^ cin;
  assign cout = (a & b) | (b & cin) | (a & cin);
endmodule
module MG_HA(
  input a,
  input b,
  output sum,
  output cout
);

  assign sum = a ^ b;
  assign cout = a & b;
endmodule
module mult16u_booth4_sklansky(
  input [15:0] multiplicand,
  input [15:0] multiplier,
  output [31:0] product
);

  wire be_2x_0_0;
  wire be_2x_0_1;
  wire be_2x_0_10;
  wire be_2x_0_11;
  wire be_2x_0_12;
  wire be_2x_0_13;
  wire be_2x_0_14;
  wire be_2x_0_15;
  wire be_2x_0_16;
  wire be_2x_0_17;
  wire be_2x_0_2;
  wire be_2x_0_3;
  wire be_2x_0_4;
  wire be_2x_0_5;
  wire be_2x_0_6;
  wire be_2x_0_7;
  wire be_2x_0_8;
  wire be_2x_0_9;
  wire be_2x_1_0;
  wire be_2x_1_1;
  wire be_2x_1_10;
  wire be_2x_1_11;
  wire be_2x_1_12;
  wire be_2x_1_13;
  wire be_2x_1_14;
  wire be_2x_1_15;
  wire be_2x_1_16;
  wire be_2x_1_17;
  wire be_2x_1_2;
  wire be_2x_1_3;
  wire be_2x_1_4;
  wire be_2x_1_5;
  wire be_2x_1_6;
  wire be_2x_1_7;
  wire be_2x_1_8;
  wire be_2x_1_9;
  wire be_2x_2_0;
  wire be_2x_2_1;
  wire be_2x_2_10;
  wire be_2x_2_11;
  wire be_2x_2_12;
  wire be_2x_2_13;
  wire be_2x_2_14;
  wire be_2x_2_15;
  wire be_2x_2_16;
  wire be_2x_2_17;
  wire be_2x_2_2;
  wire be_2x_2_3;
  wire be_2x_2_4;
  wire be_2x_2_5;
  wire be_2x_2_6;
  wire be_2x_2_7;
  wire be_2x_2_8;
  wire be_2x_2_9;
  wire be_2x_3_0;
  wire be_2x_3_1;
  wire be_2x_3_10;
  wire be_2x_3_11;
  wire be_2x_3_12;
  wire be_2x_3_13;
  wire be_2x_3_14;
  wire be_2x_3_15;
  wire be_2x_3_16;
  wire be_2x_3_17;
  wire be_2x_3_2;
  wire be_2x_3_3;
  wire be_2x_3_4;
  wire be_2x_3_5;
  wire be_2x_3_6;
  wire be_2x_3_7;
  wire be_2x_3_8;
  wire be_2x_3_9;
  wire be_2x_4_0;
  wire be_2x_4_1;
  wire be_2x_4_10;
  wire be_2x_4_11;
  wire be_2x_4_12;
  wire be_2x_4_13;
  wire be_2x_4_14;
  wire be_2x_4_15;
  wire be_2x_4_16;
  wire be_2x_4_17;
  wire be_2x_4_2;
  wire be_2x_4_3;
  wire be_2x_4_4;
  wire be_2x_4_5;
  wire be_2x_4_6;
  wire be_2x_4_7;
  wire be_2x_4_8;
  wire be_2x_4_9;
  wire be_2x_5_0;
  wire be_2x_5_1;
  wire be_2x_5_10;
  wire be_2x_5_11;
  wire be_2x_5_12;
  wire be_2x_5_13;
  wire be_2x_5_14;
  wire be_2x_5_15;
  wire be_2x_5_16;
  wire be_2x_5_17;
  wire be_2x_5_2;
  wire be_2x_5_3;
  wire be_2x_5_4;
  wire be_2x_5_5;
  wire be_2x_5_6;
  wire be_2x_5_7;
  wire be_2x_5_8;
  wire be_2x_5_9;
  wire be_2x_6_0;
  wire be_2x_6_1;
  wire be_2x_6_10;
  wire be_2x_6_11;
  wire be_2x_6_12;
  wire be_2x_6_13;
  wire be_2x_6_14;
  wire be_2x_6_15;
  wire be_2x_6_16;
  wire be_2x_6_17;
  wire be_2x_6_2;
  wire be_2x_6_3;
  wire be_2x_6_4;
  wire be_2x_6_5;
  wire be_2x_6_6;
  wire be_2x_6_7;
  wire be_2x_6_8;
  wire be_2x_6_9;
  wire be_2x_7_0;
  wire be_2x_7_1;
  wire be_2x_7_10;
  wire be_2x_7_11;
  wire be_2x_7_12;
  wire be_2x_7_13;
  wire be_2x_7_14;
  wire be_2x_7_15;
  wire be_2x_7_16;
  wire be_2x_7_17;
  wire be_2x_7_2;
  wire be_2x_7_3;
  wire be_2x_7_4;
  wire be_2x_7_5;
  wire be_2x_7_6;
  wire be_2x_7_7;
  wire be_2x_7_8;
  wire be_2x_7_9;
  wire be_2x_8_0;
  wire be_2x_8_1;
  wire be_2x_8_10;
  wire be_2x_8_11;
  wire be_2x_8_12;
  wire be_2x_8_13;
  wire be_2x_8_14;
  wire be_2x_8_15;
  wire be_2x_8_2;
  wire be_2x_8_3;
  wire be_2x_8_4;
  wire be_2x_8_5;
  wire be_2x_8_6;
  wire be_2x_8_7;
  wire be_2x_8_8;
  wire be_2x_8_9;
  wire be_c_0;
  wire be_c_1;
  wire be_c_2;
  wire be_c_3;
  wire be_c_4;
  wire be_c_5;
  wire be_c_6;
  wire be_c_7;
  wire be_c_8;
  wire be_d_0;
  wire be_d_1;
  wire be_d_2;
  wire be_d_3;
  wire be_d_4;
  wire be_d_5;
  wire be_d_6;
  wire be_d_7;
  wire be_d_8;
  wire be_neg_0;
  wire be_neg_1;
  wire be_neg_2;
  wire be_neg_3;
  wire be_neg_4;
  wire be_neg_5;
  wire be_neg_6;
  wire be_neg_7;
  wire be_neg_8;
  wire be_s1_0;
  wire be_s1_1;
  wire be_s1_2;
  wire be_s1_3;
  wire be_s1_4;
  wire be_s1_5;
  wire be_s1_6;
  wire be_s1_7;
  wire be_s1_8;
  wire be_s2_0;
  wire be_s2_1;
  wire be_s2_2;
  wire be_s2_3;
  wire be_s2_4;
  wire be_s2_5;
  wire be_s2_6;
  wire be_s2_7;
  wire be_s2_8;
  wire be_s2_a_0;
  wire be_s2_a_1;
  wire be_s2_a_2;
  wire be_s2_a_3;
  wire be_s2_a_4;
  wire be_s2_a_5;
  wire be_s2_a_6;
  wire be_s2_a_7;
  wire be_s2_a_8;
  wire be_s2_b_0;
  wire be_s2_b_1;
  wire be_s2_b_2;
  wire be_s2_b_3;
  wire be_s2_b_4;
  wire be_s2_b_5;
  wire be_s2_b_6;
  wire be_s2_b_7;
  wire be_s2_b_8;
  wire be_x_0_0;
  wire be_x_0_1;
  wire be_x_0_10;
  wire be_x_0_11;
  wire be_x_0_12;
  wire be_x_0_13;
  wire be_x_0_14;
  wire be_x_0_15;
  wire be_x_0_16;
  wire be_x_0_17;
  wire be_x_0_2;
  wire be_x_0_3;
  wire be_x_0_4;
  wire be_x_0_5;
  wire be_x_0_6;
  wire be_x_0_7;
  wire be_x_0_8;
  wire be_x_0_9;
  wire be_x_1_0;
  wire be_x_1_1;
  wire be_x_1_10;
  wire be_x_1_11;
  wire be_x_1_12;
  wire be_x_1_13;
  wire be_x_1_14;
  wire be_x_1_15;
  wire be_x_1_16;
  wire be_x_1_17;
  wire be_x_1_2;
  wire be_x_1_3;
  wire be_x_1_4;
  wire be_x_1_5;
  wire be_x_1_6;
  wire be_x_1_7;
  wire be_x_1_8;
  wire be_x_1_9;
  wire be_x_2_0;
  wire be_x_2_1;
  wire be_x_2_10;
  wire be_x_2_11;
  wire be_x_2_12;
  wire be_x_2_13;
  wire be_x_2_14;
  wire be_x_2_15;
  wire be_x_2_16;
  wire be_x_2_17;
  wire be_x_2_2;
  wire be_x_2_3;
  wire be_x_2_4;
  wire be_x_2_5;
  wire be_x_2_6;
  wire be_x_2_7;
  wire be_x_2_8;
  wire be_x_2_9;
  wire be_x_3_0;
  wire be_x_3_1;
  wire be_x_3_10;
  wire be_x_3_11;
  wire be_x_3_12;
  wire be_x_3_13;
  wire be_x_3_14;
  wire be_x_3_15;
  wire be_x_3_16;
  wire be_x_3_17;
  wire be_x_3_2;
  wire be_x_3_3;
  wire be_x_3_4;
  wire be_x_3_5;
  wire be_x_3_6;
  wire be_x_3_7;
  wire be_x_3_8;
  wire be_x_3_9;
  wire be_x_4_0;
  wire be_x_4_1;
  wire be_x_4_10;
  wire be_x_4_11;
  wire be_x_4_12;
  wire be_x_4_13;
  wire be_x_4_14;
  wire be_x_4_15;
  wire be_x_4_16;
  wire be_x_4_17;
  wire be_x_4_2;
  wire be_x_4_3;
  wire be_x_4_4;
  wire be_x_4_5;
  wire be_x_4_6;
  wire be_x_4_7;
  wire be_x_4_8;
  wire be_x_4_9;
  wire be_x_5_0;
  wire be_x_5_1;
  wire be_x_5_10;
  wire be_x_5_11;
  wire be_x_5_12;
  wire be_x_5_13;
  wire be_x_5_14;
  wire be_x_5_15;
  wire be_x_5_16;
  wire be_x_5_17;
  wire be_x_5_2;
  wire be_x_5_3;
  wire be_x_5_4;
  wire be_x_5_5;
  wire be_x_5_6;
  wire be_x_5_7;
  wire be_x_5_8;
  wire be_x_5_9;
  wire be_x_6_0;
  wire be_x_6_1;
  wire be_x_6_10;
  wire be_x_6_11;
  wire be_x_6_12;
  wire be_x_6_13;
  wire be_x_6_14;
  wire be_x_6_15;
  wire be_x_6_16;
  wire be_x_6_17;
  wire be_x_6_2;
  wire be_x_6_3;
  wire be_x_6_4;
  wire be_x_6_5;
  wire be_x_6_6;
  wire be_x_6_7;
  wire be_x_6_8;
  wire be_x_6_9;
  wire be_x_7_0;
  wire be_x_7_1;
  wire be_x_7_10;
  wire be_x_7_11;
  wire be_x_7_12;
  wire be_x_7_13;
  wire be_x_7_14;
  wire be_x_7_15;
  wire be_x_7_16;
  wire be_x_7_17;
  wire be_x_7_2;
  wire be_x_7_3;
  wire be_x_7_4;
  wire be_x_7_5;
  wire be_x_7_6;
  wire be_x_7_7;
  wire be_x_7_8;
  wire be_x_7_9;
  wire be_x_8_0;
  wire be_x_8_1;
  wire be_x_8_10;
  wire be_x_8_11;
  wire be_x_8_12;
  wire be_x_8_13;
  wire be_x_8_14;
  wire be_x_8_15;
  wire be_x_8_2;
  wire be_x_8_3;
  wire be_x_8_4;
  wire be_x_8_5;
  wire be_x_8_6;
  wire be_x_8_7;
  wire be_x_8_8;
  wire be_x_8_9;
  wire not_pp_0_19;
  wire not_pp_1_19;
  wire not_pp_2_21;
  wire not_pp_3_23;
  wire not_pp_4_25;
  wire not_pp_5_27;
  wire not_pp_6_29;
  wire not_pp_7_31;
  wire ny_0;
  wire ny_1;
  wire ny_10;
  wire ny_11;
  wire ny_12;
  wire ny_13;
  wire ny_14;
  wire ny_15;
  wire ny_2;
  wire ny_3;
  wire ny_4;
  wire ny_5;
  wire ny_6;
  wire ny_7;
  wire ny_8;
  wire ny_9;
  wire one;
  wire pp_0_0;
  wire pp_0_1;
  wire pp_0_10;
  wire pp_0_11;
  wire pp_0_12;
  wire pp_0_13;
  wire pp_0_14;
  wire pp_0_15;
  wire pp_0_16;
  wire pp_0_17;
  wire pp_0_2;
  wire pp_0_3;
  wire pp_0_4;
  wire pp_0_5;
  wire pp_0_6;
  wire pp_0_7;
  wire pp_0_8;
  wire pp_0_9;
  wire pp_1_10;
  wire pp_1_11;
  wire pp_1_12;
  wire pp_1_13;
  wire pp_1_14;
  wire pp_1_15;
  wire pp_1_16;
  wire pp_1_17;
  wire pp_1_18;
  wire pp_1_19;
  wire pp_1_2;
  wire pp_1_3;
  wire pp_1_4;
  wire pp_1_5;
  wire pp_1_6;
  wire pp_1_7;
  wire pp_1_8;
  wire pp_1_9;
  wire pp_2_10;
  wire pp_2_11;
  wire pp_2_12;
  wire pp_2_13;
  wire pp_2_14;
  wire pp_2_15;
  wire pp_2_16;
  wire pp_2_17;
  wire pp_2_18;
  wire pp_2_19;
  wire pp_2_20;
  wire pp_2_21;
  wire pp_2_4;
  wire pp_2_5;
  wire pp_2_6;
  wire pp_2_7;
  wire pp_2_8;
  wire pp_2_9;
  wire pp_3_10;
  wire pp_3_11;
  wire pp_3_12;
  wire pp_3_13;
  wire pp_3_14;
  wire pp_3_15;
  wire pp_3_16;
  wire pp_3_17;
  wire pp_3_18;
  wire pp_3_19;
  wire pp_3_20;
  wire pp_3_21;
  wire pp_3_22;
  wire pp_3_23;
  wire pp_3_6;
  wire pp_3_7;
  wire pp_3_8;
  wire pp_3_9;
  wire pp_4_10;
  wire pp_4_11;
  wire pp_4_12;
  wire pp_4_13;
  wire pp_4_14;
  wire pp_4_15;
  wire pp_4_16;
  wire pp_4_17;
  wire pp_4_18;
  wire pp_4_19;
  wire pp_4_20;
  wire pp_4_21;
  wire pp_4_22;
  wire pp_4_23;
  wire pp_4_24;
  wire pp_4_25;
  wire pp_4_8;
  wire pp_4_9;
  wire pp_5_10;
  wire pp_5_11;
  wire pp_5_12;
  wire pp_5_13;
  wire pp_5_14;
  wire pp_5_15;
  wire pp_5_16;
  wire pp_5_17;
  wire pp_5_18;
  wire pp_5_19;
  wire pp_5_20;
  wire pp_5_21;
  wire pp_5_22;
  wire pp_5_23;
  wire pp_5_24;
  wire pp_5_25;
  wire pp_5_26;
  wire pp_5_27;
  wire pp_6_12;
  wire pp_6_13;
  wire pp_6_14;
  wire pp_6_15;
  wire pp_6_16;
  wire pp_6_17;
  wire pp_6_18;
  wire pp_6_19;
  wire pp_6_20;
  wire pp_6_21;
  wire pp_6_22;
  wire pp_6_23;
  wire pp_6_24;
  wire pp_6_25;
  wire pp_6_26;
  wire pp_6_27;
  wire pp_6_28;
  wire pp_6_29;
  wire pp_7_14;
  wire pp_7_15;
  wire pp_7_16;
  wire pp_7_17;
  wire pp_7_18;
  wire pp_7_19;
  wire pp_7_20;
  wire pp_7_21;
  wire pp_7_22;
  wire pp_7_23;
  wire pp_7_24;
  wire pp_7_25;
  wire pp_7_26;
  wire pp_7_27;
  wire pp_7_28;
  wire pp_7_29;
  wire pp_7_30;
  wire pp_7_31;
  wire pp_8_16;
  wire pp_8_17;
  wire pp_8_18;
  wire pp_8_19;
  wire pp_8_20;
  wire pp_8_21;
  wire pp_8_22;
  wire pp_8_23;
  wire pp_8_24;
  wire pp_8_25;
  wire pp_8_26;
  wire pp_8_27;
  wire pp_8_28;
  wire pp_8_29;
  wire pp_8_30;
  wire pp_8_31;
  wire px_0_0;
  wire px_0_1;
  wire px_0_10;
  wire px_0_11;
  wire px_0_12;
  wire px_0_13;
  wire px_0_14;
  wire px_0_15;
  wire px_0_16;
  wire px_0_17;
  wire px_0_18;
  wire px_0_2;
  wire px_0_3;
  wire px_0_4;
  wire px_0_5;
  wire px_0_6;
  wire px_0_7;
  wire px_0_8;
  wire px_0_9;
  wire px_1_0;
  wire px_1_1;
  wire px_1_10;
  wire px_1_11;
  wire px_1_12;
  wire px_1_13;
  wire px_1_14;
  wire px_1_15;
  wire px_1_16;
  wire px_1_17;
  wire px_1_18;
  wire px_1_2;
  wire px_1_3;
  wire px_1_4;
  wire px_1_5;
  wire px_1_6;
  wire px_1_7;
  wire px_1_8;
  wire px_1_9;
  wire px_2_0;
  wire px_2_1;
  wire px_2_10;
  wire px_2_11;
  wire px_2_12;
  wire px_2_13;
  wire px_2_14;
  wire px_2_15;
  wire px_2_16;
  wire px_2_17;
  wire px_2_18;
  wire px_2_2;
  wire px_2_3;
  wire px_2_4;
  wire px_2_5;
  wire px_2_6;
  wire px_2_7;
  wire px_2_8;
  wire px_2_9;
  wire px_3_0;
  wire px_3_1;
  wire px_3_10;
  wire px_3_11;
  wire px_3_12;
  wire px_3_13;
  wire px_3_14;
  wire px_3_15;
  wire px_3_16;
  wire px_3_17;
  wire px_3_18;
  wire px_3_2;
  wire px_3_3;
  wire px_3_4;
  wire px_3_5;
  wire px_3_6;
  wire px_3_7;
  wire px_3_8;
  wire px_3_9;
  wire px_4_0;
  wire px_4_1;
  wire px_4_10;
  wire px_4_11;
  wire px_4_12;
  wire px_4_13;
  wire px_4_14;
  wire px_4_15;
  wire px_4_16;
  wire px_4_17;
  wire px_4_18;
  wire px_4_2;
  wire px_4_3;
  wire px_4_4;
  wire px_4_5;
  wire px_4_6;
  wire px_4_7;
  wire px_4_8;
  wire px_4_9;
  wire px_5_0;
  wire px_5_1;
  wire px_5_10;
  wire px_5_11;
  wire px_5_12;
  wire px_5_13;
  wire px_5_14;
  wire px_5_15;
  wire px_5_16;
  wire px_5_17;
  wire px_5_18;
  wire px_5_2;
  wire px_5_3;
  wire px_5_4;
  wire px_5_5;
  wire px_5_6;
  wire px_5_7;
  wire px_5_8;
  wire px_5_9;
  wire px_6_0;
  wire px_6_1;
  wire px_6_10;
  wire px_6_11;
  wire px_6_12;
  wire px_6_13;
  wire px_6_14;
  wire px_6_15;
  wire px_6_16;
  wire px_6_17;
  wire px_6_18;
  wire px_6_2;
  wire px_6_3;
  wire px_6_4;
  wire px_6_5;
  wire px_6_6;
  wire px_6_7;
  wire px_6_8;
  wire px_6_9;
  wire px_7_0;
  wire px_7_1;
  wire px_7_10;
  wire px_7_11;
  wire px_7_12;
  wire px_7_13;
  wire px_7_14;
  wire px_7_15;
  wire px_7_16;
  wire px_7_17;
  wire px_7_18;
  wire px_7_2;
  wire px_7_3;
  wire px_7_4;
  wire px_7_5;
  wire px_7_6;
  wire px_7_7;
  wire px_7_8;
  wire px_7_9;
  wire px_8_0;
  wire px_8_1;
  wire px_8_10;
  wire px_8_11;
  wire px_8_12;
  wire px_8_13;
  wire px_8_14;
  wire px_8_15;
  wire px_8_16;
  wire px_8_17;
  wire px_8_18;
  wire px_8_2;
  wire px_8_3;
  wire px_8_4;
  wire px_8_5;
  wire px_8_6;
  wire px_8_7;
  wire px_8_8;
  wire px_8_9;
  wire x_0;
  wire x_1;
  wire x_10;
  wire x_11;
  wire x_12;
  wire x_13;
  wire x_14;
  wire x_15;
  wire x_2;
  wire x_3;
  wire x_4;
  wire x_5;
  wire x_6;
  wire x_7;
  wire x_8;
  wire x_9;
  wire y_0;
  wire y_1;
  wire y_10;
  wire y_11;
  wire y_12;
  wire y_13;
  wire y_14;
  wire y_15;
  wire y_2;
  wire y_3;
  wire y_4;
  wire y_5;
  wire y_6;
  wire y_7;
  wire y_8;
  wire y_9;
  wire zero;
  assign be_2x_0_0 = ~(px_0_0 & be_s2_0);
  assign be_2x_0_1 = ~(px_0_1 & be_s2_0);
  assign be_2x_0_10 = ~(px_0_10 & be_s2_0);
  assign be_2x_0_11 = ~(px_0_11 & be_s2_0);
  assign be_2x_0_12 = ~(px_0_12 & be_s2_0);
  assign be_2x_0_13 = ~(px_0_13 & be_s2_0);
  assign be_2x_0_14 = ~(px_0_14 & be_s2_0);
  assign be_2x_0_15 = ~(px_0_15 & be_s2_0);
  assign be_2x_0_16 = ~(px_0_16 & be_s2_0);
  assign be_2x_0_17 = ~(px_0_17 & be_s2_0);
  assign be_2x_0_2 = ~(px_0_2 & be_s2_0);
  assign be_2x_0_3 = ~(px_0_3 & be_s2_0);
  assign be_2x_0_4 = ~(px_0_4 & be_s2_0);
  assign be_2x_0_5 = ~(px_0_5 & be_s2_0);
  assign be_2x_0_6 = ~(px_0_6 & be_s2_0);
  assign be_2x_0_7 = ~(px_0_7 & be_s2_0);
  assign be_2x_0_8 = ~(px_0_8 & be_s2_0);
  assign be_2x_0_9 = ~(px_0_9 & be_s2_0);
  assign be_2x_1_0 = ~(px_1_0 & be_s2_1);
  assign be_2x_1_1 = ~(px_1_1 & be_s2_1);
  assign be_2x_1_10 = ~(px_1_10 & be_s2_1);
  assign be_2x_1_11 = ~(px_1_11 & be_s2_1);
  assign be_2x_1_12 = ~(px_1_12 & be_s2_1);
  assign be_2x_1_13 = ~(px_1_13 & be_s2_1);
  assign be_2x_1_14 = ~(px_1_14 & be_s2_1);
  assign be_2x_1_15 = ~(px_1_15 & be_s2_1);
  assign be_2x_1_16 = ~(px_1_16 & be_s2_1);
  assign be_2x_1_17 = ~(px_1_17 & be_s2_1);
  assign be_2x_1_2 = ~(px_1_2 & be_s2_1);
  assign be_2x_1_3 = ~(px_1_3 & be_s2_1);
  assign be_2x_1_4 = ~(px_1_4 & be_s2_1);
  assign be_2x_1_5 = ~(px_1_5 & be_s2_1);
  assign be_2x_1_6 = ~(px_1_6 & be_s2_1);
  assign be_2x_1_7 = ~(px_1_7 & be_s2_1);
  assign be_2x_1_8 = ~(px_1_8 & be_s2_1);
  assign be_2x_1_9 = ~(px_1_9 & be_s2_1);
  assign be_2x_2_0 = ~(px_2_0 & be_s2_2);
  assign be_2x_2_1 = ~(px_2_1 & be_s2_2);
  assign be_2x_2_10 = ~(px_2_10 & be_s2_2);
  assign be_2x_2_11 = ~(px_2_11 & be_s2_2);
  assign be_2x_2_12 = ~(px_2_12 & be_s2_2);
  assign be_2x_2_13 = ~(px_2_13 & be_s2_2);
  assign be_2x_2_14 = ~(px_2_14 & be_s2_2);
  assign be_2x_2_15 = ~(px_2_15 & be_s2_2);
  assign be_2x_2_16 = ~(px_2_16 & be_s2_2);
  assign be_2x_2_17 = ~(px_2_17 & be_s2_2);
  assign be_2x_2_2 = ~(px_2_2 & be_s2_2);
  assign be_2x_2_3 = ~(px_2_3 & be_s2_2);
  assign be_2x_2_4 = ~(px_2_4 & be_s2_2);
  assign be_2x_2_5 = ~(px_2_5 & be_s2_2);
  assign be_2x_2_6 = ~(px_2_6 & be_s2_2);
  assign be_2x_2_7 = ~(px_2_7 & be_s2_2);
  assign be_2x_2_8 = ~(px_2_8 & be_s2_2);
  assign be_2x_2_9 = ~(px_2_9 & be_s2_2);
  assign be_2x_3_0 = ~(px_3_0 & be_s2_3);
  assign be_2x_3_1 = ~(px_3_1 & be_s2_3);
  assign be_2x_3_10 = ~(px_3_10 & be_s2_3);
  assign be_2x_3_11 = ~(px_3_11 & be_s2_3);
  assign be_2x_3_12 = ~(px_3_12 & be_s2_3);
  assign be_2x_3_13 = ~(px_3_13 & be_s2_3);
  assign be_2x_3_14 = ~(px_3_14 & be_s2_3);
  assign be_2x_3_15 = ~(px_3_15 & be_s2_3);
  assign be_2x_3_16 = ~(px_3_16 & be_s2_3);
  assign be_2x_3_17 = ~(px_3_17 & be_s2_3);
  assign be_2x_3_2 = ~(px_3_2 & be_s2_3);
  assign be_2x_3_3 = ~(px_3_3 & be_s2_3);
  assign be_2x_3_4 = ~(px_3_4 & be_s2_3);
  assign be_2x_3_5 = ~(px_3_5 & be_s2_3);
  assign be_2x_3_6 = ~(px_3_6 & be_s2_3);
  assign be_2x_3_7 = ~(px_3_7 & be_s2_3);
  assign be_2x_3_8 = ~(px_3_8 & be_s2_3);
  assign be_2x_3_9 = ~(px_3_9 & be_s2_3);
  assign be_2x_4_0 = ~(px_4_0 & be_s2_4);
  assign be_2x_4_1 = ~(px_4_1 & be_s2_4);
  assign be_2x_4_10 = ~(px_4_10 & be_s2_4);
  assign be_2x_4_11 = ~(px_4_11 & be_s2_4);
  assign be_2x_4_12 = ~(px_4_12 & be_s2_4);
  assign be_2x_4_13 = ~(px_4_13 & be_s2_4);
  assign be_2x_4_14 = ~(px_4_14 & be_s2_4);
  assign be_2x_4_15 = ~(px_4_15 & be_s2_4);
  assign be_2x_4_16 = ~(px_4_16 & be_s2_4);
  assign be_2x_4_17 = ~(px_4_17 & be_s2_4);
  assign be_2x_4_2 = ~(px_4_2 & be_s2_4);
  assign be_2x_4_3 = ~(px_4_3 & be_s2_4);
  assign be_2x_4_4 = ~(px_4_4 & be_s2_4);
  assign be_2x_4_5 = ~(px_4_5 & be_s2_4);
  assign be_2x_4_6 = ~(px_4_6 & be_s2_4);
  assign be_2x_4_7 = ~(px_4_7 & be_s2_4);
  assign be_2x_4_8 = ~(px_4_8 & be_s2_4);
  assign be_2x_4_9 = ~(px_4_9 & be_s2_4);
  assign be_2x_5_0 = ~(px_5_0 & be_s2_5);
  assign be_2x_5_1 = ~(px_5_1 & be_s2_5);
  assign be_2x_5_10 = ~(px_5_10 & be_s2_5);
  assign be_2x_5_11 = ~(px_5_11 & be_s2_5);
  assign be_2x_5_12 = ~(px_5_12 & be_s2_5);
  assign be_2x_5_13 = ~(px_5_13 & be_s2_5);
  assign be_2x_5_14 = ~(px_5_14 & be_s2_5);
  assign be_2x_5_15 = ~(px_5_15 & be_s2_5);
  assign be_2x_5_16 = ~(px_5_16 & be_s2_5);
  assign be_2x_5_17 = ~(px_5_17 & be_s2_5);
  assign be_2x_5_2 = ~(px_5_2 & be_s2_5);
  assign be_2x_5_3 = ~(px_5_3 & be_s2_5);
  assign be_2x_5_4 = ~(px_5_4 & be_s2_5);
  assign be_2x_5_5 = ~(px_5_5 & be_s2_5);
  assign be_2x_5_6 = ~(px_5_6 & be_s2_5);
  assign be_2x_5_7 = ~(px_5_7 & be_s2_5);
  assign be_2x_5_8 = ~(px_5_8 & be_s2_5);
  assign be_2x_5_9 = ~(px_5_9 & be_s2_5);
  assign be_2x_6_0 = ~(px_6_0 & be_s2_6);
  assign be_2x_6_1 = ~(px_6_1 & be_s2_6);
  assign be_2x_6_10 = ~(px_6_10 & be_s2_6);
  assign be_2x_6_11 = ~(px_6_11 & be_s2_6);
  assign be_2x_6_12 = ~(px_6_12 & be_s2_6);
  assign be_2x_6_13 = ~(px_6_13 & be_s2_6);
  assign be_2x_6_14 = ~(px_6_14 & be_s2_6);
  assign be_2x_6_15 = ~(px_6_15 & be_s2_6);
  assign be_2x_6_16 = ~(px_6_16 & be_s2_6);
  assign be_2x_6_17 = ~(px_6_17 & be_s2_6);
  assign be_2x_6_2 = ~(px_6_2 & be_s2_6);
  assign be_2x_6_3 = ~(px_6_3 & be_s2_6);
  assign be_2x_6_4 = ~(px_6_4 & be_s2_6);
  assign be_2x_6_5 = ~(px_6_5 & be_s2_6);
  assign be_2x_6_6 = ~(px_6_6 & be_s2_6);
  assign be_2x_6_7 = ~(px_6_7 & be_s2_6);
  assign be_2x_6_8 = ~(px_6_8 & be_s2_6);
  assign be_2x_6_9 = ~(px_6_9 & be_s2_6);
  assign be_2x_7_0 = ~(px_7_0 & be_s2_7);
  assign be_2x_7_1 = ~(px_7_1 & be_s2_7);
  assign be_2x_7_10 = ~(px_7_10 & be_s2_7);
  assign be_2x_7_11 = ~(px_7_11 & be_s2_7);
  assign be_2x_7_12 = ~(px_7_12 & be_s2_7);
  assign be_2x_7_13 = ~(px_7_13 & be_s2_7);
  assign be_2x_7_14 = ~(px_7_14 & be_s2_7);
  assign be_2x_7_15 = ~(px_7_15 & be_s2_7);
  assign be_2x_7_16 = ~(px_7_16 & be_s2_7);
  assign be_2x_7_17 = ~(px_7_17 & be_s2_7);
  assign be_2x_7_2 = ~(px_7_2 & be_s2_7);
  assign be_2x_7_3 = ~(px_7_3 & be_s2_7);
  assign be_2x_7_4 = ~(px_7_4 & be_s2_7);
  assign be_2x_7_5 = ~(px_7_5 & be_s2_7);
  assign be_2x_7_6 = ~(px_7_6 & be_s2_7);
  assign be_2x_7_7 = ~(px_7_7 & be_s2_7);
  assign be_2x_7_8 = ~(px_7_8 & be_s2_7);
  assign be_2x_7_9 = ~(px_7_9 & be_s2_7);
  assign be_2x_8_0 = ~(px_8_0 & be_s2_8);
  assign be_2x_8_1 = ~(px_8_1 & be_s2_8);
  assign be_2x_8_10 = ~(px_8_10 & be_s2_8);
  assign be_2x_8_11 = ~(px_8_11 & be_s2_8);
  assign be_2x_8_12 = ~(px_8_12 & be_s2_8);
  assign be_2x_8_13 = ~(px_8_13 & be_s2_8);
  assign be_2x_8_14 = ~(px_8_14 & be_s2_8);
  assign be_2x_8_15 = ~(px_8_15 & be_s2_8);
  assign be_2x_8_2 = ~(px_8_2 & be_s2_8);
  assign be_2x_8_3 = ~(px_8_3 & be_s2_8);
  assign be_2x_8_4 = ~(px_8_4 & be_s2_8);
  assign be_2x_8_5 = ~(px_8_5 & be_s2_8);
  assign be_2x_8_6 = ~(px_8_6 & be_s2_8);
  assign be_2x_8_7 = ~(px_8_7 & be_s2_8);
  assign be_2x_8_8 = ~(px_8_8 & be_s2_8);
  assign be_2x_8_9 = ~(px_8_9 & be_s2_8);
  assign be_c_0 = be_d_0 & be_neg_0;
  assign be_c_1 = be_d_1 & be_neg_1;
  assign be_c_2 = be_d_2 & be_neg_2;
  assign be_c_3 = be_d_3 & be_neg_3;
  assign be_c_4 = be_d_4 & be_neg_4;
  assign be_c_5 = be_d_5 & be_neg_5;
  assign be_c_6 = be_d_6 & be_neg_6;
  assign be_c_7 = be_d_7 & be_neg_7;
  assign be_c_8 = be_d_8 & be_neg_8;
  assign be_d_0 = ny_0 | one;
  assign be_d_1 = ny_2 | ny_1;
  assign be_d_2 = ny_4 | ny_3;
  assign be_d_3 = ny_6 | ny_5;
  assign be_d_4 = ny_8 | ny_7;
  assign be_d_5 = ny_10 | ny_9;
  assign be_d_6 = ny_12 | ny_11;
  assign be_d_7 = ny_14 | ny_13;
  assign be_d_8 = one | ny_15;
  assign be_neg_0 = y_1;
  assign be_neg_1 = y_3;
  assign be_neg_2 = y_5;
  assign be_neg_3 = y_7;
  assign be_neg_4 = y_9;
  assign be_neg_5 = y_11;
  assign be_neg_6 = y_13;
  assign be_neg_7 = y_15;
  assign be_neg_8 = zero;
  assign be_s1_0 = y_0 ^ zero;
  assign be_s1_1 = y_2 ^ y_1;
  assign be_s1_2 = y_4 ^ y_3;
  assign be_s1_3 = y_6 ^ y_5;
  assign be_s1_4 = y_8 ^ y_7;
  assign be_s1_5 = y_10 ^ y_9;
  assign be_s1_6 = y_12 ^ y_11;
  assign be_s1_7 = y_14 ^ y_13;
  assign be_s1_8 = zero ^ y_15;
  assign be_s2_0 = be_s2_a_0 | be_s2_b_0;
  assign be_s2_1 = be_s2_a_1 | be_s2_b_1;
  assign be_s2_2 = be_s2_a_2 | be_s2_b_2;
  assign be_s2_3 = be_s2_a_3 | be_s2_b_3;
  assign be_s2_4 = be_s2_a_4 | be_s2_b_4;
  assign be_s2_5 = be_s2_a_5 | be_s2_b_5;
  assign be_s2_6 = be_s2_a_6 | be_s2_b_6;
  assign be_s2_7 = be_s2_a_7 | be_s2_b_7;
  assign be_s2_8 = be_s2_a_8 | be_s2_b_8;
  assign be_s2_a_0 = ny_1 & y_0 & zero;
  assign be_s2_a_1 = ny_3 & y_2 & y_1;
  assign be_s2_a_2 = ny_5 & y_4 & y_3;
  assign be_s2_a_3 = ny_7 & y_6 & y_5;
  assign be_s2_a_4 = ny_9 & y_8 & y_7;
  assign be_s2_a_5 = ny_11 & y_10 & y_9;
  assign be_s2_a_6 = ny_13 & y_12 & y_11;
  assign be_s2_a_7 = ny_15 & y_14 & y_13;
  assign be_s2_a_8 = one & zero & y_15;
  assign be_s2_b_0 = y_1 & ny_0 & one;
  assign be_s2_b_1 = y_3 & ny_2 & ny_1;
  assign be_s2_b_2 = y_5 & ny_4 & ny_3;
  assign be_s2_b_3 = y_7 & ny_6 & ny_5;
  assign be_s2_b_4 = y_9 & ny_8 & ny_7;
  assign be_s2_b_5 = y_11 & ny_10 & ny_9;
  assign be_s2_b_6 = y_13 & ny_12 & ny_11;
  assign be_s2_b_7 = y_15 & ny_14 & ny_13;
  assign be_s2_b_8 = zero & one & ny_15;
  assign be_x_0_0 = ~(px_0_1 & be_s1_0);
  assign be_x_0_1 = ~(px_0_2 & be_s1_0);
  assign be_x_0_10 = ~(px_0_11 & be_s1_0);
  assign be_x_0_11 = ~(px_0_12 & be_s1_0);
  assign be_x_0_12 = ~(px_0_13 & be_s1_0);
  assign be_x_0_13 = ~(px_0_14 & be_s1_0);
  assign be_x_0_14 = ~(px_0_15 & be_s1_0);
  assign be_x_0_15 = ~(px_0_16 & be_s1_0);
  assign be_x_0_16 = ~(px_0_17 & be_s1_0);
  assign be_x_0_17 = ~(px_0_18 & be_s1_0);
  assign be_x_0_2 = ~(px_0_3 & be_s1_0);
  assign be_x_0_3 = ~(px_0_4 & be_s1_0);
  assign be_x_0_4 = ~(px_0_5 & be_s1_0);
  assign be_x_0_5 = ~(px_0_6 & be_s1_0);
  assign be_x_0_6 = ~(px_0_7 & be_s1_0);
  assign be_x_0_7 = ~(px_0_8 & be_s1_0);
  assign be_x_0_8 = ~(px_0_9 & be_s1_0);
  assign be_x_0_9 = ~(px_0_10 & be_s1_0);
  assign be_x_1_0 = ~(px_1_1 & be_s1_1);
  assign be_x_1_1 = ~(px_1_2 & be_s1_1);
  assign be_x_1_10 = ~(px_1_11 & be_s1_1);
  assign be_x_1_11 = ~(px_1_12 & be_s1_1);
  assign be_x_1_12 = ~(px_1_13 & be_s1_1);
  assign be_x_1_13 = ~(px_1_14 & be_s1_1);
  assign be_x_1_14 = ~(px_1_15 & be_s1_1);
  assign be_x_1_15 = ~(px_1_16 & be_s1_1);
  assign be_x_1_16 = ~(px_1_17 & be_s1_1);
  assign be_x_1_17 = ~(px_1_18 & be_s1_1);
  assign be_x_1_2 = ~(px_1_3 & be_s1_1);
  assign be_x_1_3 = ~(px_1_4 & be_s1_1);
  assign be_x_1_4 = ~(px_1_5 & be_s1_1);
  assign be_x_1_5 = ~(px_1_6 & be_s1_1);
  assign be_x_1_6 = ~(px_1_7 & be_s1_1);
  assign be_x_1_7 = ~(px_1_8 & be_s1_1);
  assign be_x_1_8 = ~(px_1_9 & be_s1_1);
  assign be_x_1_9 = ~(px_1_10 & be_s1_1);
  assign be_x_2_0 = ~(px_2_1 & be_s1_2);
  assign be_x_2_1 = ~(px_2_2 & be_s1_2);
  assign be_x_2_10 = ~(px_2_11 & be_s1_2);
  assign be_x_2_11 = ~(px_2_12 & be_s1_2);
  assign be_x_2_12 = ~(px_2_13 & be_s1_2);
  assign be_x_2_13 = ~(px_2_14 & be_s1_2);
  assign be_x_2_14 = ~(px_2_15 & be_s1_2);
  assign be_x_2_15 = ~(px_2_16 & be_s1_2);
  assign be_x_2_16 = ~(px_2_17 & be_s1_2);
  assign be_x_2_17 = ~(px_2_18 & be_s1_2);
  assign be_x_2_2 = ~(px_2_3 & be_s1_2);
  assign be_x_2_3 = ~(px_2_4 & be_s1_2);
  assign be_x_2_4 = ~(px_2_5 & be_s1_2);
  assign be_x_2_5 = ~(px_2_6 & be_s1_2);
  assign be_x_2_6 = ~(px_2_7 & be_s1_2);
  assign be_x_2_7 = ~(px_2_8 & be_s1_2);
  assign be_x_2_8 = ~(px_2_9 & be_s1_2);
  assign be_x_2_9 = ~(px_2_10 & be_s1_2);
  assign be_x_3_0 = ~(px_3_1 & be_s1_3);
  assign be_x_3_1 = ~(px_3_2 & be_s1_3);
  assign be_x_3_10 = ~(px_3_11 & be_s1_3);
  assign be_x_3_11 = ~(px_3_12 & be_s1_3);
  assign be_x_3_12 = ~(px_3_13 & be_s1_3);
  assign be_x_3_13 = ~(px_3_14 & be_s1_3);
  assign be_x_3_14 = ~(px_3_15 & be_s1_3);
  assign be_x_3_15 = ~(px_3_16 & be_s1_3);
  assign be_x_3_16 = ~(px_3_17 & be_s1_3);
  assign be_x_3_17 = ~(px_3_18 & be_s1_3);
  assign be_x_3_2 = ~(px_3_3 & be_s1_3);
  assign be_x_3_3 = ~(px_3_4 & be_s1_3);
  assign be_x_3_4 = ~(px_3_5 & be_s1_3);
  assign be_x_3_5 = ~(px_3_6 & be_s1_3);
  assign be_x_3_6 = ~(px_3_7 & be_s1_3);
  assign be_x_3_7 = ~(px_3_8 & be_s1_3);
  assign be_x_3_8 = ~(px_3_9 & be_s1_3);
  assign be_x_3_9 = ~(px_3_10 & be_s1_3);
  assign be_x_4_0 = ~(px_4_1 & be_s1_4);
  assign be_x_4_1 = ~(px_4_2 & be_s1_4);
  assign be_x_4_10 = ~(px_4_11 & be_s1_4);
  assign be_x_4_11 = ~(px_4_12 & be_s1_4);
  assign be_x_4_12 = ~(px_4_13 & be_s1_4);
  assign be_x_4_13 = ~(px_4_14 & be_s1_4);
  assign be_x_4_14 = ~(px_4_15 & be_s1_4);
  assign be_x_4_15 = ~(px_4_16 & be_s1_4);
  assign be_x_4_16 = ~(px_4_17 & be_s1_4);
  assign be_x_4_17 = ~(px_4_18 & be_s1_4);
  assign be_x_4_2 = ~(px_4_3 & be_s1_4);
  assign be_x_4_3 = ~(px_4_4 & be_s1_4);
  assign be_x_4_4 = ~(px_4_5 & be_s1_4);
  assign be_x_4_5 = ~(px_4_6 & be_s1_4);
  assign be_x_4_6 = ~(px_4_7 & be_s1_4);
  assign be_x_4_7 = ~(px_4_8 & be_s1_4);
  assign be_x_4_8 = ~(px_4_9 & be_s1_4);
  assign be_x_4_9 = ~(px_4_10 & be_s1_4);
  assign be_x_5_0 = ~(px_5_1 & be_s1_5);
  assign be_x_5_1 = ~(px_5_2 & be_s1_5);
  assign be_x_5_10 = ~(px_5_11 & be_s1_5);
  assign be_x_5_11 = ~(px_5_12 & be_s1_5);
  assign be_x_5_12 = ~(px_5_13 & be_s1_5);
  assign be_x_5_13 = ~(px_5_14 & be_s1_5);
  assign be_x_5_14 = ~(px_5_15 & be_s1_5);
  assign be_x_5_15 = ~(px_5_16 & be_s1_5);
  assign be_x_5_16 = ~(px_5_17 & be_s1_5);
  assign be_x_5_17 = ~(px_5_18 & be_s1_5);
  assign be_x_5_2 = ~(px_5_3 & be_s1_5);
  assign be_x_5_3 = ~(px_5_4 & be_s1_5);
  assign be_x_5_4 = ~(px_5_5 & be_s1_5);
  assign be_x_5_5 = ~(px_5_6 & be_s1_5);
  assign be_x_5_6 = ~(px_5_7 & be_s1_5);
  assign be_x_5_7 = ~(px_5_8 & be_s1_5);
  assign be_x_5_8 = ~(px_5_9 & be_s1_5);
  assign be_x_5_9 = ~(px_5_10 & be_s1_5);
  assign be_x_6_0 = ~(px_6_1 & be_s1_6);
  assign be_x_6_1 = ~(px_6_2 & be_s1_6);
  assign be_x_6_10 = ~(px_6_11 & be_s1_6);
  assign be_x_6_11 = ~(px_6_12 & be_s1_6);
  assign be_x_6_12 = ~(px_6_13 & be_s1_6);
  assign be_x_6_13 = ~(px_6_14 & be_s1_6);
  assign be_x_6_14 = ~(px_6_15 & be_s1_6);
  assign be_x_6_15 = ~(px_6_16 & be_s1_6);
  assign be_x_6_16 = ~(px_6_17 & be_s1_6);
  assign be_x_6_17 = ~(px_6_18 & be_s1_6);
  assign be_x_6_2 = ~(px_6_3 & be_s1_6);
  assign be_x_6_3 = ~(px_6_4 & be_s1_6);
  assign be_x_6_4 = ~(px_6_5 & be_s1_6);
  assign be_x_6_5 = ~(px_6_6 & be_s1_6);
  assign be_x_6_6 = ~(px_6_7 & be_s1_6);
  assign be_x_6_7 = ~(px_6_8 & be_s1_6);
  assign be_x_6_8 = ~(px_6_9 & be_s1_6);
  assign be_x_6_9 = ~(px_6_10 & be_s1_6);
  assign be_x_7_0 = ~(px_7_1 & be_s1_7);
  assign be_x_7_1 = ~(px_7_2 & be_s1_7);
  assign be_x_7_10 = ~(px_7_11 & be_s1_7);
  assign be_x_7_11 = ~(px_7_12 & be_s1_7);
  assign be_x_7_12 = ~(px_7_13 & be_s1_7);
  assign be_x_7_13 = ~(px_7_14 & be_s1_7);
  assign be_x_7_14 = ~(px_7_15 & be_s1_7);
  assign be_x_7_15 = ~(px_7_16 & be_s1_7);
  assign be_x_7_16 = ~(px_7_17 & be_s1_7);
  assign be_x_7_17 = ~(px_7_18 & be_s1_7);
  assign be_x_7_2 = ~(px_7_3 & be_s1_7);
  assign be_x_7_3 = ~(px_7_4 & be_s1_7);
  assign be_x_7_4 = ~(px_7_5 & be_s1_7);
  assign be_x_7_5 = ~(px_7_6 & be_s1_7);
  assign be_x_7_6 = ~(px_7_7 & be_s1_7);
  assign be_x_7_7 = ~(px_7_8 & be_s1_7);
  assign be_x_7_8 = ~(px_7_9 & be_s1_7);
  assign be_x_7_9 = ~(px_7_10 & be_s1_7);
  assign be_x_8_0 = ~(px_8_1 & be_s1_8);
  assign be_x_8_1 = ~(px_8_2 & be_s1_8);
  assign be_x_8_10 = ~(px_8_11 & be_s1_8);
  assign be_x_8_11 = ~(px_8_12 & be_s1_8);
  assign be_x_8_12 = ~(px_8_13 & be_s1_8);
  assign be_x_8_13 = ~(px_8_14 & be_s1_8);
  assign be_x_8_14 = ~(px_8_15 & be_s1_8);
  assign be_x_8_15 = ~(px_8_16 & be_s1_8);
  assign be_x_8_2 = ~(px_8_3 & be_s1_8);
  assign be_x_8_3 = ~(px_8_4 & be_s1_8);
  assign be_x_8_4 = ~(px_8_5 & be_s1_8);
  assign be_x_8_5 = ~(px_8_6 & be_s1_8);
  assign be_x_8_6 = ~(px_8_7 & be_s1_8);
  assign be_x_8_7 = ~(px_8_8 & be_s1_8);
  assign be_x_8_8 = ~(px_8_9 & be_s1_8);
  assign be_x_8_9 = ~(px_8_10 & be_s1_8);
  assign not_pp_0_19 = ~pp_0_17;
  assign not_pp_1_19 = ~pp_1_19;
  assign not_pp_2_21 = ~pp_2_21;
  assign not_pp_3_23 = ~pp_3_23;
  assign not_pp_4_25 = ~pp_4_25;
  assign not_pp_5_27 = ~pp_5_27;
  assign not_pp_6_29 = ~pp_6_29;
  assign not_pp_7_31 = ~pp_7_31;
  assign ny_0 = ~multiplier[0];
  assign ny_1 = ~multiplier[1];
  assign ny_10 = ~multiplier[10];
  assign ny_11 = ~multiplier[11];
  assign ny_12 = ~multiplier[12];
  assign ny_13 = ~multiplier[13];
  assign ny_14 = ~multiplier[14];
  assign ny_15 = ~multiplier[15];
  assign ny_2 = ~multiplier[2];
  assign ny_3 = ~multiplier[3];
  assign ny_4 = ~multiplier[4];
  assign ny_5 = ~multiplier[5];
  assign ny_6 = ~multiplier[6];
  assign ny_7 = ~multiplier[7];
  assign ny_8 = ~multiplier[8];
  assign ny_9 = ~multiplier[9];
  assign one = 1'b1;
  assign pp_0_0 = ~(be_2x_0_0 & be_x_0_0);
  assign pp_0_1 = ~(be_2x_0_1 & be_x_0_1);
  assign pp_0_10 = ~(be_2x_0_10 & be_x_0_10);
  assign pp_0_11 = ~(be_2x_0_11 & be_x_0_11);
  assign pp_0_12 = ~(be_2x_0_12 & be_x_0_12);
  assign pp_0_13 = ~(be_2x_0_13 & be_x_0_13);
  assign pp_0_14 = ~(be_2x_0_14 & be_x_0_14);
  assign pp_0_15 = ~(be_2x_0_15 & be_x_0_15);
  assign pp_0_16 = ~(be_2x_0_16 & be_x_0_16);
  assign pp_0_17 = ~(be_2x_0_17 & be_x_0_17);
  assign pp_0_2 = ~(be_2x_0_2 & be_x_0_2);
  assign pp_0_3 = ~(be_2x_0_3 & be_x_0_3);
  assign pp_0_4 = ~(be_2x_0_4 & be_x_0_4);
  assign pp_0_5 = ~(be_2x_0_5 & be_x_0_5);
  assign pp_0_6 = ~(be_2x_0_6 & be_x_0_6);
  assign pp_0_7 = ~(be_2x_0_7 & be_x_0_7);
  assign pp_0_8 = ~(be_2x_0_8 & be_x_0_8);
  assign pp_0_9 = ~(be_2x_0_9 & be_x_0_9);
  assign pp_1_10 = ~(be_2x_1_8 & be_x_1_8);
  assign pp_1_11 = ~(be_2x_1_9 & be_x_1_9);
  assign pp_1_12 = ~(be_2x_1_10 & be_x_1_10);
  assign pp_1_13 = ~(be_2x_1_11 & be_x_1_11);
  assign pp_1_14 = ~(be_2x_1_12 & be_x_1_12);
  assign pp_1_15 = ~(be_2x_1_13 & be_x_1_13);
  assign pp_1_16 = ~(be_2x_1_14 & be_x_1_14);
  assign pp_1_17 = ~(be_2x_1_15 & be_x_1_15);
  assign pp_1_18 = ~(be_2x_1_16 & be_x_1_16);
  assign pp_1_19 = ~(be_2x_1_17 & be_x_1_17);
  assign pp_1_2 = ~(be_2x_1_0 & be_x_1_0);
  assign pp_1_3 = ~(be_2x_1_1 & be_x_1_1);
  assign pp_1_4 = ~(be_2x_1_2 & be_x_1_2);
  assign pp_1_5 = ~(be_2x_1_3 & be_x_1_3);
  assign pp_1_6 = ~(be_2x_1_4 & be_x_1_4);
  assign pp_1_7 = ~(be_2x_1_5 & be_x_1_5);
  assign pp_1_8 = ~(be_2x_1_6 & be_x_1_6);
  assign pp_1_9 = ~(be_2x_1_7 & be_x_1_7);
  assign pp_2_10 = ~(be_2x_2_6 & be_x_2_6);
  assign pp_2_11 = ~(be_2x_2_7 & be_x_2_7);
  assign pp_2_12 = ~(be_2x_2_8 & be_x_2_8);
  assign pp_2_13 = ~(be_2x_2_9 & be_x_2_9);
  assign pp_2_14 = ~(be_2x_2_10 & be_x_2_10);
  assign pp_2_15 = ~(be_2x_2_11 & be_x_2_11);
  assign pp_2_16 = ~(be_2x_2_12 & be_x_2_12);
  assign pp_2_17 = ~(be_2x_2_13 & be_x_2_13);
  assign pp_2_18 = ~(be_2x_2_14 & be_x_2_14);
  assign pp_2_19 = ~(be_2x_2_15 & be_x_2_15);
  assign pp_2_20 = ~(be_2x_2_16 & be_x_2_16);
  assign pp_2_21 = ~(be_2x_2_17 & be_x_2_17);
  assign pp_2_4 = ~(be_2x_2_0 & be_x_2_0);
  assign pp_2_5 = ~(be_2x_2_1 & be_x_2_1);
  assign pp_2_6 = ~(be_2x_2_2 & be_x_2_2);
  assign pp_2_7 = ~(be_2x_2_3 & be_x_2_3);
  assign pp_2_8 = ~(be_2x_2_4 & be_x_2_4);
  assign pp_2_9 = ~(be_2x_2_5 & be_x_2_5);
  assign pp_3_10 = ~(be_2x_3_4 & be_x_3_4);
  assign pp_3_11 = ~(be_2x_3_5 & be_x_3_5);
  assign pp_3_12 = ~(be_2x_3_6 & be_x_3_6);
  assign pp_3_13 = ~(be_2x_3_7 & be_x_3_7);
  assign pp_3_14 = ~(be_2x_3_8 & be_x_3_8);
  assign pp_3_15 = ~(be_2x_3_9 & be_x_3_9);
  assign pp_3_16 = ~(be_2x_3_10 & be_x_3_10);
  assign pp_3_17 = ~(be_2x_3_11 & be_x_3_11);
  assign pp_3_18 = ~(be_2x_3_12 & be_x_3_12);
  assign pp_3_19 = ~(be_2x_3_13 & be_x_3_13);
  assign pp_3_20 = ~(be_2x_3_14 & be_x_3_14);
  assign pp_3_21 = ~(be_2x_3_15 & be_x_3_15);
  assign pp_3_22 = ~(be_2x_3_16 & be_x_3_16);
  assign pp_3_23 = ~(be_2x_3_17 & be_x_3_17);
  assign pp_3_6 = ~(be_2x_3_0 & be_x_3_0);
  assign pp_3_7 = ~(be_2x_3_1 & be_x_3_1);
  assign pp_3_8 = ~(be_2x_3_2 & be_x_3_2);
  assign pp_3_9 = ~(be_2x_3_3 & be_x_3_3);
  assign pp_4_10 = ~(be_2x_4_2 & be_x_4_2);
  assign pp_4_11 = ~(be_2x_4_3 & be_x_4_3);
  assign pp_4_12 = ~(be_2x_4_4 & be_x_4_4);
  assign pp_4_13 = ~(be_2x_4_5 & be_x_4_5);
  assign pp_4_14 = ~(be_2x_4_6 & be_x_4_6);
  assign pp_4_15 = ~(be_2x_4_7 & be_x_4_7);
  assign pp_4_16 = ~(be_2x_4_8 & be_x_4_8);
  assign pp_4_17 = ~(be_2x_4_9 & be_x_4_9);
  assign pp_4_18 = ~(be_2x_4_10 & be_x_4_10);
  assign pp_4_19 = ~(be_2x_4_11 & be_x_4_11);
  assign pp_4_20 = ~(be_2x_4_12 & be_x_4_12);
  assign pp_4_21 = ~(be_2x_4_13 & be_x_4_13);
  assign pp_4_22 = ~(be_2x_4_14 & be_x_4_14);
  assign pp_4_23 = ~(be_2x_4_15 & be_x_4_15);
  assign pp_4_24 = ~(be_2x_4_16 & be_x_4_16);
  assign pp_4_25 = ~(be_2x_4_17 & be_x_4_17);
  assign pp_4_8 = ~(be_2x_4_0 & be_x_4_0);
  assign pp_4_9 = ~(be_2x_4_1 & be_x_4_1);
  assign pp_5_10 = ~(be_2x_5_0 & be_x_5_0);
  assign pp_5_11 = ~(be_2x_5_1 & be_x_5_1);
  assign pp_5_12 = ~(be_2x_5_2 & be_x_5_2);
  assign pp_5_13 = ~(be_2x_5_3 & be_x_5_3);
  assign pp_5_14 = ~(be_2x_5_4 & be_x_5_4);
  assign pp_5_15 = ~(be_2x_5_5 & be_x_5_5);
  assign pp_5_16 = ~(be_2x_5_6 & be_x_5_6);
  assign pp_5_17 = ~(be_2x_5_7 & be_x_5_7);
  assign pp_5_18 = ~(be_2x_5_8 & be_x_5_8);
  assign pp_5_19 = ~(be_2x_5_9 & be_x_5_9);
  assign pp_5_20 = ~(be_2x_5_10 & be_x_5_10);
  assign pp_5_21 = ~(be_2x_5_11 & be_x_5_11);
  assign pp_5_22 = ~(be_2x_5_12 & be_x_5_12);
  assign pp_5_23 = ~(be_2x_5_13 & be_x_5_13);
  assign pp_5_24 = ~(be_2x_5_14 & be_x_5_14);
  assign pp_5_25 = ~(be_2x_5_15 & be_x_5_15);
  assign pp_5_26 = ~(be_2x_5_16 & be_x_5_16);
  assign pp_5_27 = ~(be_2x_5_17 & be_x_5_17);
  assign pp_6_12 = ~(be_2x_6_0 & be_x_6_0);
  assign pp_6_13 = ~(be_2x_6_1 & be_x_6_1);
  assign pp_6_14 = ~(be_2x_6_2 & be_x_6_2);
  assign pp_6_15 = ~(be_2x_6_3 & be_x_6_3);
  assign pp_6_16 = ~(be_2x_6_4 & be_x_6_4);
  assign pp_6_17 = ~(be_2x_6_5 & be_x_6_5);
  assign pp_6_18 = ~(be_2x_6_6 & be_x_6_6);
  assign pp_6_19 = ~(be_2x_6_7 & be_x_6_7);
  assign pp_6_20 = ~(be_2x_6_8 & be_x_6_8);
  assign pp_6_21 = ~(be_2x_6_9 & be_x_6_9);
  assign pp_6_22 = ~(be_2x_6_10 & be_x_6_10);
  assign pp_6_23 = ~(be_2x_6_11 & be_x_6_11);
  assign pp_6_24 = ~(be_2x_6_12 & be_x_6_12);
  assign pp_6_25 = ~(be_2x_6_13 & be_x_6_13);
  assign pp_6_26 = ~(be_2x_6_14 & be_x_6_14);
  assign pp_6_27 = ~(be_2x_6_15 & be_x_6_15);
  assign pp_6_28 = ~(be_2x_6_16 & be_x_6_16);
  assign pp_6_29 = ~(be_2x_6_17 & be_x_6_17);
  assign pp_7_14 = ~(be_2x_7_0 & be_x_7_0);
  assign pp_7_15 = ~(be_2x_7_1 & be_x_7_1);
  assign pp_7_16 = ~(be_2x_7_2 & be_x_7_2);
  assign pp_7_17 = ~(be_2x_7_3 & be_x_7_3);
  assign pp_7_18 = ~(be_2x_7_4 & be_x_7_4);
  assign pp_7_19 = ~(be_2x_7_5 & be_x_7_5);
  assign pp_7_20 = ~(be_2x_7_6 & be_x_7_6);
  assign pp_7_21 = ~(be_2x_7_7 & be_x_7_7);
  assign pp_7_22 = ~(be_2x_7_8 & be_x_7_8);
  assign pp_7_23 = ~(be_2x_7_9 & be_x_7_9);
  assign pp_7_24 = ~(be_2x_7_10 & be_x_7_10);
  assign pp_7_25 = ~(be_2x_7_11 & be_x_7_11);
  assign pp_7_26 = ~(be_2x_7_12 & be_x_7_12);
  assign pp_7_27 = ~(be_2x_7_13 & be_x_7_13);
  assign pp_7_28 = ~(be_2x_7_14 & be_x_7_14);
  assign pp_7_29 = ~(be_2x_7_15 & be_x_7_15);
  assign pp_7_30 = ~(be_2x_7_16 & be_x_7_16);
  assign pp_7_31 = ~(be_2x_7_17 & be_x_7_17);
  assign pp_8_16 = ~(be_2x_8_0 & be_x_8_0);
  assign pp_8_17 = ~(be_2x_8_1 & be_x_8_1);
  assign pp_8_18 = ~(be_2x_8_2 & be_x_8_2);
  assign pp_8_19 = ~(be_2x_8_3 & be_x_8_3);
  assign pp_8_20 = ~(be_2x_8_4 & be_x_8_4);
  assign pp_8_21 = ~(be_2x_8_5 & be_x_8_5);
  assign pp_8_22 = ~(be_2x_8_6 & be_x_8_6);
  assign pp_8_23 = ~(be_2x_8_7 & be_x_8_7);
  assign pp_8_24 = ~(be_2x_8_8 & be_x_8_8);
  assign pp_8_25 = ~(be_2x_8_9 & be_x_8_9);
  assign pp_8_26 = ~(be_2x_8_10 & be_x_8_10);
  assign pp_8_27 = ~(be_2x_8_11 & be_x_8_11);
  assign pp_8_28 = ~(be_2x_8_12 & be_x_8_12);
  assign pp_8_29 = ~(be_2x_8_13 & be_x_8_13);
  assign pp_8_30 = ~(be_2x_8_14 & be_x_8_14);
  assign pp_8_31 = ~(be_2x_8_15 & be_x_8_15);
  assign px_0_0 = be_neg_0;
  assign px_0_1 = be_neg_0 ^ x_0;
  assign px_0_10 = be_neg_0 ^ x_9;
  assign px_0_11 = be_neg_0 ^ x_10;
  assign px_0_12 = be_neg_0 ^ x_11;
  assign px_0_13 = be_neg_0 ^ x_12;
  assign px_0_14 = be_neg_0 ^ x_13;
  assign px_0_15 = be_neg_0 ^ x_14;
  assign px_0_16 = be_neg_0 ^ x_15;
  assign px_0_17 = be_neg_0 ^ zero;
  assign px_0_18 = be_neg_0 ^ zero;
  assign px_0_2 = be_neg_0 ^ x_1;
  assign px_0_3 = be_neg_0 ^ x_2;
  assign px_0_4 = be_neg_0 ^ x_3;
  assign px_0_5 = be_neg_0 ^ x_4;
  assign px_0_6 = be_neg_0 ^ x_5;
  assign px_0_7 = be_neg_0 ^ x_6;
  assign px_0_8 = be_neg_0 ^ x_7;
  assign px_0_9 = be_neg_0 ^ x_8;
  assign px_1_0 = be_neg_1;
  assign px_1_1 = be_neg_1 ^ x_0;
  assign px_1_10 = be_neg_1 ^ x_9;
  assign px_1_11 = be_neg_1 ^ x_10;
  assign px_1_12 = be_neg_1 ^ x_11;
  assign px_1_13 = be_neg_1 ^ x_12;
  assign px_1_14 = be_neg_1 ^ x_13;
  assign px_1_15 = be_neg_1 ^ x_14;
  assign px_1_16 = be_neg_1 ^ x_15;
  assign px_1_17 = be_neg_1 ^ zero;
  assign px_1_18 = be_neg_1 ^ zero;
  assign px_1_2 = be_neg_1 ^ x_1;
  assign px_1_3 = be_neg_1 ^ x_2;
  assign px_1_4 = be_neg_1 ^ x_3;
  assign px_1_5 = be_neg_1 ^ x_4;
  assign px_1_6 = be_neg_1 ^ x_5;
  assign px_1_7 = be_neg_1 ^ x_6;
  assign px_1_8 = be_neg_1 ^ x_7;
  assign px_1_9 = be_neg_1 ^ x_8;
  assign px_2_0 = be_neg_2;
  assign px_2_1 = be_neg_2 ^ x_0;
  assign px_2_10 = be_neg_2 ^ x_9;
  assign px_2_11 = be_neg_2 ^ x_10;
  assign px_2_12 = be_neg_2 ^ x_11;
  assign px_2_13 = be_neg_2 ^ x_12;
  assign px_2_14 = be_neg_2 ^ x_13;
  assign px_2_15 = be_neg_2 ^ x_14;
  assign px_2_16 = be_neg_2 ^ x_15;
  assign px_2_17 = be_neg_2 ^ zero;
  assign px_2_18 = be_neg_2 ^ zero;
  assign px_2_2 = be_neg_2 ^ x_1;
  assign px_2_3 = be_neg_2 ^ x_2;
  assign px_2_4 = be_neg_2 ^ x_3;
  assign px_2_5 = be_neg_2 ^ x_4;
  assign px_2_6 = be_neg_2 ^ x_5;
  assign px_2_7 = be_neg_2 ^ x_6;
  assign px_2_8 = be_neg_2 ^ x_7;
  assign px_2_9 = be_neg_2 ^ x_8;
  assign px_3_0 = be_neg_3;
  assign px_3_1 = be_neg_3 ^ x_0;
  assign px_3_10 = be_neg_3 ^ x_9;
  assign px_3_11 = be_neg_3 ^ x_10;
  assign px_3_12 = be_neg_3 ^ x_11;
  assign px_3_13 = be_neg_3 ^ x_12;
  assign px_3_14 = be_neg_3 ^ x_13;
  assign px_3_15 = be_neg_3 ^ x_14;
  assign px_3_16 = be_neg_3 ^ x_15;
  assign px_3_17 = be_neg_3 ^ zero;
  assign px_3_18 = be_neg_3 ^ zero;
  assign px_3_2 = be_neg_3 ^ x_1;
  assign px_3_3 = be_neg_3 ^ x_2;
  assign px_3_4 = be_neg_3 ^ x_3;
  assign px_3_5 = be_neg_3 ^ x_4;
  assign px_3_6 = be_neg_3 ^ x_5;
  assign px_3_7 = be_neg_3 ^ x_6;
  assign px_3_8 = be_neg_3 ^ x_7;
  assign px_3_9 = be_neg_3 ^ x_8;
  assign px_4_0 = be_neg_4;
  assign px_4_1 = be_neg_4 ^ x_0;
  assign px_4_10 = be_neg_4 ^ x_9;
  assign px_4_11 = be_neg_4 ^ x_10;
  assign px_4_12 = be_neg_4 ^ x_11;
  assign px_4_13 = be_neg_4 ^ x_12;
  assign px_4_14 = be_neg_4 ^ x_13;
  assign px_4_15 = be_neg_4 ^ x_14;
  assign px_4_16 = be_neg_4 ^ x_15;
  assign px_4_17 = be_neg_4 ^ zero;
  assign px_4_18 = be_neg_4 ^ zero;
  assign px_4_2 = be_neg_4 ^ x_1;
  assign px_4_3 = be_neg_4 ^ x_2;
  assign px_4_4 = be_neg_4 ^ x_3;
  assign px_4_5 = be_neg_4 ^ x_4;
  assign px_4_6 = be_neg_4 ^ x_5;
  assign px_4_7 = be_neg_4 ^ x_6;
  assign px_4_8 = be_neg_4 ^ x_7;
  assign px_4_9 = be_neg_4 ^ x_8;
  assign px_5_0 = be_neg_5;
  assign px_5_1 = be_neg_5 ^ x_0;
  assign px_5_10 = be_neg_5 ^ x_9;
  assign px_5_11 = be_neg_5 ^ x_10;
  assign px_5_12 = be_neg_5 ^ x_11;
  assign px_5_13 = be_neg_5 ^ x_12;
  assign px_5_14 = be_neg_5 ^ x_13;
  assign px_5_15 = be_neg_5 ^ x_14;
  assign px_5_16 = be_neg_5 ^ x_15;
  assign px_5_17 = be_neg_5 ^ zero;
  assign px_5_18 = be_neg_5 ^ zero;
  assign px_5_2 = be_neg_5 ^ x_1;
  assign px_5_3 = be_neg_5 ^ x_2;
  assign px_5_4 = be_neg_5 ^ x_3;
  assign px_5_5 = be_neg_5 ^ x_4;
  assign px_5_6 = be_neg_5 ^ x_5;
  assign px_5_7 = be_neg_5 ^ x_6;
  assign px_5_8 = be_neg_5 ^ x_7;
  assign px_5_9 = be_neg_5 ^ x_8;
  assign px_6_0 = be_neg_6;
  assign px_6_1 = be_neg_6 ^ x_0;
  assign px_6_10 = be_neg_6 ^ x_9;
  assign px_6_11 = be_neg_6 ^ x_10;
  assign px_6_12 = be_neg_6 ^ x_11;
  assign px_6_13 = be_neg_6 ^ x_12;
  assign px_6_14 = be_neg_6 ^ x_13;
  assign px_6_15 = be_neg_6 ^ x_14;
  assign px_6_16 = be_neg_6 ^ x_15;
  assign px_6_17 = be_neg_6 ^ zero;
  assign px_6_18 = be_neg_6 ^ zero;
  assign px_6_2 = be_neg_6 ^ x_1;
  assign px_6_3 = be_neg_6 ^ x_2;
  assign px_6_4 = be_neg_6 ^ x_3;
  assign px_6_5 = be_neg_6 ^ x_4;
  assign px_6_6 = be_neg_6 ^ x_5;
  assign px_6_7 = be_neg_6 ^ x_6;
  assign px_6_8 = be_neg_6 ^ x_7;
  assign px_6_9 = be_neg_6 ^ x_8;
  assign px_7_0 = be_neg_7;
  assign px_7_1 = be_neg_7 ^ x_0;
  assign px_7_10 = be_neg_7 ^ x_9;
  assign px_7_11 = be_neg_7 ^ x_10;
  assign px_7_12 = be_neg_7 ^ x_11;
  assign px_7_13 = be_neg_7 ^ x_12;
  assign px_7_14 = be_neg_7 ^ x_13;
  assign px_7_15 = be_neg_7 ^ x_14;
  assign px_7_16 = be_neg_7 ^ x_15;
  assign px_7_17 = be_neg_7 ^ zero;
  assign px_7_18 = be_neg_7 ^ zero;
  assign px_7_2 = be_neg_7 ^ x_1;
  assign px_7_3 = be_neg_7 ^ x_2;
  assign px_7_4 = be_neg_7 ^ x_3;
  assign px_7_5 = be_neg_7 ^ x_4;
  assign px_7_6 = be_neg_7 ^ x_5;
  assign px_7_7 = be_neg_7 ^ x_6;
  assign px_7_8 = be_neg_7 ^ x_7;
  assign px_7_9 = be_neg_7 ^ x_8;
  assign px_8_0 = be_neg_8;
  assign px_8_1 = be_neg_8 ^ x_0;
  assign px_8_10 = be_neg_8 ^ x_9;
  assign px_8_11 = be_neg_8 ^ x_10;
  assign px_8_12 = be_neg_8 ^ x_11;
  assign px_8_13 = be_neg_8 ^ x_12;
  assign px_8_14 = be_neg_8 ^ x_13;
  assign px_8_15 = be_neg_8 ^ x_14;
  assign px_8_16 = be_neg_8 ^ x_15;
  assign px_8_17 = be_neg_8 ^ zero;
  assign px_8_18 = be_neg_8 ^ zero;
  assign px_8_2 = be_neg_8 ^ x_1;
  assign px_8_3 = be_neg_8 ^ x_2;
  assign px_8_4 = be_neg_8 ^ x_3;
  assign px_8_5 = be_neg_8 ^ x_4;
  assign px_8_6 = be_neg_8 ^ x_5;
  assign px_8_7 = be_neg_8 ^ x_6;
  assign px_8_8 = be_neg_8 ^ x_7;
  assign px_8_9 = be_neg_8 ^ x_8;
  assign x_0 = multiplicand[0];
  assign x_1 = multiplicand[1];
  assign x_10 = multiplicand[10];
  assign x_11 = multiplicand[11];
  assign x_12 = multiplicand[12];
  assign x_13 = multiplicand[13];
  assign x_14 = multiplicand[14];
  assign x_15 = multiplicand[15];
  assign x_2 = multiplicand[2];
  assign x_3 = multiplicand[3];
  assign x_4 = multiplicand[4];
  assign x_5 = multiplicand[5];
  assign x_6 = multiplicand[6];
  assign x_7 = multiplicand[7];
  assign x_8 = multiplicand[8];
  assign x_9 = multiplicand[9];
  assign y_0 = multiplier[0];
  assign y_1 = multiplier[1];
  assign y_10 = multiplier[10];
  assign y_11 = multiplier[11];
  assign y_12 = multiplier[12];
  assign y_13 = multiplier[13];
  assign y_14 = multiplier[14];
  assign y_15 = multiplier[15];
  assign y_2 = multiplier[2];
  assign y_3 = multiplier[3];
  assign y_4 = multiplier[4];
  assign y_5 = multiplier[5];
  assign y_6 = multiplier[6];
  assign y_7 = multiplier[7];
  assign y_8 = multiplier[8];
  assign y_9 = multiplier[9];
  assign zero = 1'b0;
  wire pp_0_0_0;
  wire pp_0_0_1;
  wire pp_0_1_0;
  wire pp_0_2_0;
  wire pp_0_2_1;
  wire pp_0_2_2;
  wire pp_0_3_0;
  wire pp_0_3_1;
  wire pp_0_4_0;
  wire pp_0_4_1;
  wire pp_0_4_2;
  wire pp_0_4_3;
  wire pp_0_5_0;
  wire pp_0_5_1;
  wire pp_0_5_2;
  wire pp_0_6_0;
  wire pp_0_6_1;
  wire pp_0_6_2;
  wire pp_0_6_3;
  wire pp_0_6_4;
  wire pp_0_7_0;
  wire pp_0_7_1;
  wire pp_0_7_2;
  wire pp_0_7_3;
  wire pp_0_8_0;
  wire pp_0_8_1;
  wire pp_0_8_2;
  wire pp_0_8_3;
  wire pp_0_8_4;
  wire pp_0_8_5;
  wire pp_0_9_0;
  wire pp_0_9_1;
  wire pp_0_9_2;
  wire pp_0_9_3;
  wire pp_0_9_4;
  wire pp_0_10_0;
  wire pp_0_10_1;
  wire pp_0_10_2;
  wire pp_0_10_3;
  wire pp_0_10_4;
  wire pp_0_10_5;
  wire pp_0_10_6;
  wire pp_0_11_0;
  wire pp_0_11_1;
  wire pp_0_11_2;
  wire pp_0_11_3;
  wire pp_0_11_4;
  wire pp_0_11_5;
  wire pp_0_12_0;
  wire pp_0_12_1;
  wire pp_0_12_2;
  wire pp_0_12_3;
  wire pp_0_12_4;
  wire pp_0_12_5;
  wire pp_0_12_6;
  wire pp_0_12_7;
  wire pp_0_13_0;
  wire pp_0_13_1;
  wire pp_0_13_2;
  wire pp_0_13_3;
  wire pp_0_13_4;
  wire pp_0_13_5;
  wire pp_0_13_6;
  wire pp_0_14_0;
  wire pp_0_14_1;
  wire pp_0_14_2;
  wire pp_0_14_3;
  wire pp_0_14_4;
  wire pp_0_14_5;
  wire pp_0_14_6;
  wire pp_0_14_7;
  wire pp_0_14_8;
  wire pp_0_15_0;
  wire pp_0_15_1;
  wire pp_0_15_2;
  wire pp_0_15_3;
  wire pp_0_15_4;
  wire pp_0_15_5;
  wire pp_0_15_6;
  wire pp_0_15_7;
  wire pp_0_16_0;
  wire pp_0_16_1;
  wire pp_0_16_2;
  wire pp_0_16_3;
  wire pp_0_16_4;
  wire pp_0_16_5;
  wire pp_0_16_6;
  wire pp_0_16_7;
  wire pp_0_16_8;
  wire pp_0_17_0;
  wire pp_0_17_1;
  wire pp_0_17_2;
  wire pp_0_17_3;
  wire pp_0_17_4;
  wire pp_0_17_5;
  wire pp_0_17_6;
  wire pp_0_17_7;
  wire pp_0_17_8;
  wire pp_0_18_0;
  wire pp_0_18_1;
  wire pp_0_18_2;
  wire pp_0_18_3;
  wire pp_0_18_4;
  wire pp_0_18_5;
  wire pp_0_18_6;
  wire pp_0_18_7;
  wire pp_0_18_8;
  wire pp_0_19_0;
  wire pp_0_19_1;
  wire pp_0_19_2;
  wire pp_0_19_3;
  wire pp_0_19_4;
  wire pp_0_19_5;
  wire pp_0_19_6;
  wire pp_0_19_7;
  wire pp_0_19_8;
  wire pp_0_20_0;
  wire pp_0_20_1;
  wire pp_0_20_2;
  wire pp_0_20_3;
  wire pp_0_20_4;
  wire pp_0_20_5;
  wire pp_0_20_6;
  wire pp_0_20_7;
  wire pp_0_21_0;
  wire pp_0_21_1;
  wire pp_0_21_2;
  wire pp_0_21_3;
  wire pp_0_21_4;
  wire pp_0_21_5;
  wire pp_0_21_6;
  wire pp_0_22_0;
  wire pp_0_22_1;
  wire pp_0_22_2;
  wire pp_0_22_3;
  wire pp_0_22_4;
  wire pp_0_22_5;
  wire pp_0_22_6;
  wire pp_0_23_0;
  wire pp_0_23_1;
  wire pp_0_23_2;
  wire pp_0_23_3;
  wire pp_0_23_4;
  wire pp_0_23_5;
  wire pp_0_24_0;
  wire pp_0_24_1;
  wire pp_0_24_2;
  wire pp_0_24_3;
  wire pp_0_24_4;
  wire pp_0_24_5;
  wire pp_0_25_0;
  wire pp_0_25_1;
  wire pp_0_25_2;
  wire pp_0_25_3;
  wire pp_0_25_4;
  wire pp_0_26_0;
  wire pp_0_26_1;
  wire pp_0_26_2;
  wire pp_0_26_3;
  wire pp_0_26_4;
  wire pp_0_27_0;
  wire pp_0_27_1;
  wire pp_0_27_2;
  wire pp_0_27_3;
  wire pp_0_28_0;
  wire pp_0_28_1;
  wire pp_0_28_2;
  wire pp_0_28_3;
  wire pp_0_29_0;
  wire pp_0_29_1;
  wire pp_0_29_2;
  wire pp_0_30_0;
  wire pp_0_30_1;
  wire pp_0_30_2;
  wire pp_0_31_0;
  wire pp_0_31_1;
  wire pp_1_0_0;
  wire pp_1_0_1;
  wire pp_1_1_0;
  wire pp_1_2_0;
  wire pp_1_2_1;
  wire pp_1_2_2;
  wire pp_1_3_0;
  wire pp_1_4_0;
  wire pp_1_4_1;
  wire pp_1_4_2;
  wire pp_1_4_3;
  wire pp_1_4_4;
  wire pp_1_5_0;
  wire pp_1_6_0;
  wire pp_1_6_1;
  wire pp_1_6_2;
  wire pp_1_7_0;
  wire pp_1_7_1;
  wire pp_1_7_2;
  wire pp_1_7_3;
  wire pp_1_8_0;
  wire pp_1_8_1;
  wire pp_1_8_2;
  wire pp_1_9_0;
  wire pp_1_9_1;
  wire pp_1_9_2;
  wire pp_1_9_3;
  wire pp_1_9_4;
  wire pp_1_10_0;
  wire pp_1_10_1;
  wire pp_1_10_2;
  wire pp_1_10_3;
  wire pp_1_11_0;
  wire pp_1_11_1;
  wire pp_1_11_2;
  wire pp_1_11_3;
  wire pp_1_11_4;
  wire pp_1_11_5;
  wire pp_1_12_0;
  wire pp_1_12_1;
  wire pp_1_12_2;
  wire pp_1_12_3;
  wire pp_1_13_0;
  wire pp_1_13_1;
  wire pp_1_13_2;
  wire pp_1_13_3;
  wire pp_1_13_4;
  wire pp_1_13_5;
  wire pp_1_14_0;
  wire pp_1_14_1;
  wire pp_1_14_2;
  wire pp_1_14_3;
  wire pp_1_14_4;
  wire pp_1_14_5;
  wire pp_1_15_0;
  wire pp_1_15_1;
  wire pp_1_15_2;
  wire pp_1_15_3;
  wire pp_1_15_4;
  wire pp_1_15_5;
  wire pp_1_16_0;
  wire pp_1_16_1;
  wire pp_1_16_2;
  wire pp_1_16_3;
  wire pp_1_16_4;
  wire pp_1_16_5;
  wire pp_1_17_0;
  wire pp_1_17_1;
  wire pp_1_17_2;
  wire pp_1_17_3;
  wire pp_1_17_4;
  wire pp_1_17_5;
  wire pp_1_18_0;
  wire pp_1_18_1;
  wire pp_1_18_2;
  wire pp_1_18_3;
  wire pp_1_18_4;
  wire pp_1_18_5;
  wire pp_1_19_0;
  wire pp_1_19_1;
  wire pp_1_19_2;
  wire pp_1_19_3;
  wire pp_1_19_4;
  wire pp_1_19_5;
  wire pp_1_20_0;
  wire pp_1_20_1;
  wire pp_1_20_2;
  wire pp_1_20_3;
  wire pp_1_20_4;
  wire pp_1_20_5;
  wire pp_1_21_0;
  wire pp_1_21_1;
  wire pp_1_21_2;
  wire pp_1_21_3;
  wire pp_1_21_4;
  wire pp_1_21_5;
  wire pp_1_22_0;
  wire pp_1_22_1;
  wire pp_1_22_2;
  wire pp_1_22_3;
  wire pp_1_22_4;
  wire pp_1_22_5;
  wire pp_1_23_0;
  wire pp_1_23_1;
  wire pp_1_23_2;
  wire pp_1_23_3;
  wire pp_1_24_0;
  wire pp_1_24_1;
  wire pp_1_24_2;
  wire pp_1_24_3;
  wire pp_1_24_4;
  wire pp_1_24_5;
  wire pp_1_25_0;
  wire pp_1_25_1;
  wire pp_1_25_2;
  wire pp_1_25_3;
  wire pp_1_25_4;
  wire pp_1_25_5;
  wire pp_1_26_0;
  wire pp_1_26_1;
  wire pp_1_26_2;
  wire pp_1_27_0;
  wire pp_1_27_1;
  wire pp_1_27_2;
  wire pp_1_28_0;
  wire pp_1_28_1;
  wire pp_1_28_2;
  wire pp_1_29_0;
  wire pp_1_29_1;
  wire pp_1_29_2;
  wire pp_1_29_3;
  wire pp_1_30_0;
  wire pp_1_30_1;
  wire pp_1_30_2;
  wire pp_1_31_0;
  wire pp_1_31_1;
  wire pp_2_0_0;
  wire pp_2_0_1;
  wire pp_2_1_0;
  wire pp_2_2_0;
  wire pp_2_2_1;
  wire pp_2_2_2;
  wire pp_2_3_0;
  wire pp_2_4_0;
  wire pp_2_4_1;
  wire pp_2_4_2;
  wire pp_2_5_0;
  wire pp_2_5_1;
  wire pp_2_6_0;
  wire pp_2_7_0;
  wire pp_2_7_1;
  wire pp_2_7_2;
  wire pp_2_8_0;
  wire pp_2_8_1;
  wire pp_2_9_0;
  wire pp_2_9_1;
  wire pp_2_9_2;
  wire pp_2_9_3;
  wire pp_2_10_0;
  wire pp_2_10_1;
  wire pp_2_10_2;
  wire pp_2_11_0;
  wire pp_2_11_1;
  wire pp_2_11_2;
  wire pp_2_12_0;
  wire pp_2_12_1;
  wire pp_2_12_2;
  wire pp_2_12_3;
  wire pp_2_12_4;
  wire pp_2_12_5;
  wire pp_2_13_0;
  wire pp_2_13_1;
  wire pp_2_14_0;
  wire pp_2_14_1;
  wire pp_2_14_2;
  wire pp_2_14_3;
  wire pp_2_15_0;
  wire pp_2_15_1;
  wire pp_2_15_2;
  wire pp_2_15_3;
  wire pp_2_15_4;
  wire pp_2_15_5;
  wire pp_2_16_0;
  wire pp_2_16_1;
  wire pp_2_16_2;
  wire pp_2_17_0;
  wire pp_2_17_1;
  wire pp_2_17_2;
  wire pp_2_17_3;
  wire pp_2_18_0;
  wire pp_2_18_1;
  wire pp_2_18_2;
  wire pp_2_18_3;
  wire pp_2_18_4;
  wire pp_2_18_5;
  wire pp_2_19_0;
  wire pp_2_19_1;
  wire pp_2_19_2;
  wire pp_2_20_0;
  wire pp_2_20_1;
  wire pp_2_20_2;
  wire pp_2_20_3;
  wire pp_2_21_0;
  wire pp_2_21_1;
  wire pp_2_21_2;
  wire pp_2_21_3;
  wire pp_2_22_0;
  wire pp_2_22_1;
  wire pp_2_22_2;
  wire pp_2_22_3;
  wire pp_2_23_0;
  wire pp_2_23_1;
  wire pp_2_23_2;
  wire pp_2_23_3;
  wire pp_2_24_0;
  wire pp_2_24_1;
  wire pp_2_24_2;
  wire pp_2_24_3;
  wire pp_2_24_4;
  wire pp_2_24_5;
  wire pp_2_25_0;
  wire pp_2_25_1;
  wire pp_2_25_2;
  wire pp_2_26_0;
  wire pp_2_26_1;
  wire pp_2_26_2;
  wire pp_2_27_0;
  wire pp_2_27_1;
  wire pp_2_28_0;
  wire pp_2_28_1;
  wire pp_2_29_0;
  wire pp_2_29_1;
  wire pp_2_29_2;
  wire pp_2_30_0;
  wire pp_2_30_1;
  wire pp_2_31_0;
  wire pp_2_31_1;
  wire pp_2_31_2;
  wire pp_3_0_0;
  wire pp_3_0_1;
  wire pp_3_1_0;
  wire pp_3_2_0;
  wire pp_3_2_1;
  wire pp_3_3_0;
  wire pp_3_3_1;
  wire pp_3_4_0;
  wire pp_3_4_1;
  wire pp_3_5_0;
  wire pp_3_5_1;
  wire pp_3_5_2;
  wire pp_3_6_0;
  wire pp_3_7_0;
  wire pp_3_7_1;
  wire pp_3_8_0;
  wire pp_3_8_1;
  wire pp_3_9_0;
  wire pp_3_9_1;
  wire pp_3_9_2;
  wire pp_3_10_0;
  wire pp_3_10_1;
  wire pp_3_10_2;
  wire pp_3_11_0;
  wire pp_3_11_1;
  wire pp_3_11_2;
  wire pp_3_12_0;
  wire pp_3_12_1;
  wire pp_3_12_2;
  wire pp_3_13_0;
  wire pp_3_13_1;
  wire pp_3_13_2;
  wire pp_3_14_0;
  wire pp_3_14_1;
  wire pp_3_14_2;
  wire pp_3_15_0;
  wire pp_3_15_1;
  wire pp_3_15_2;
  wire pp_3_16_0;
  wire pp_3_16_1;
  wire pp_3_16_2;
  wire pp_3_17_0;
  wire pp_3_17_1;
  wire pp_3_17_2;
  wire pp_3_18_0;
  wire pp_3_18_1;
  wire pp_3_18_2;
  wire pp_3_19_0;
  wire pp_3_19_1;
  wire pp_3_19_2;
  wire pp_3_20_0;
  wire pp_3_20_1;
  wire pp_3_20_2;
  wire pp_3_21_0;
  wire pp_3_21_1;
  wire pp_3_21_2;
  wire pp_3_22_0;
  wire pp_3_22_1;
  wire pp_3_22_2;
  wire pp_3_23_0;
  wire pp_3_23_1;
  wire pp_3_23_2;
  wire pp_3_24_0;
  wire pp_3_24_1;
  wire pp_3_24_2;
  wire pp_3_25_0;
  wire pp_3_25_1;
  wire pp_3_25_2;
  wire pp_3_26_0;
  wire pp_3_26_1;
  wire pp_3_26_2;
  wire pp_3_27_0;
  wire pp_3_27_1;
  wire pp_3_27_2;
  wire pp_3_28_0;
  wire pp_3_29_0;
  wire pp_3_29_1;
  wire pp_3_30_0;
  wire pp_3_30_1;
  wire pp_3_30_2;
  wire pp_3_31_0;
  wire pp_4_0_0;
  wire pp_4_0_1;
  wire pp_4_1_0;
  wire pp_4_2_0;
  wire pp_4_2_1;
  wire pp_4_3_0;
  wire pp_4_3_1;
  wire pp_4_4_0;
  wire pp_4_4_1;
  wire pp_4_5_0;
  wire pp_4_5_1;
  wire pp_4_6_0;
  wire pp_4_6_1;
  wire pp_4_7_0;
  wire pp_4_7_1;
  wire pp_4_8_0;
  wire pp_4_8_1;
  wire pp_4_9_0;
  wire pp_4_9_1;
  wire pp_4_10_0;
  wire pp_4_10_1;
  wire pp_4_11_0;
  wire pp_4_11_1;
  wire pp_4_12_0;
  wire pp_4_12_1;
  wire pp_4_13_0;
  wire pp_4_13_1;
  wire pp_4_14_0;
  wire pp_4_14_1;
  wire pp_4_15_0;
  wire pp_4_15_1;
  wire pp_4_16_0;
  wire pp_4_16_1;
  wire pp_4_17_0;
  wire pp_4_17_1;
  wire pp_4_18_0;
  wire pp_4_18_1;
  wire pp_4_19_0;
  wire pp_4_19_1;
  wire pp_4_20_0;
  wire pp_4_20_1;
  wire pp_4_21_0;
  wire pp_4_21_1;
  wire pp_4_22_0;
  wire pp_4_22_1;
  wire pp_4_23_0;
  wire pp_4_23_1;
  wire pp_4_24_0;
  wire pp_4_24_1;
  wire pp_4_25_0;
  wire pp_4_25_1;
  wire pp_4_26_0;
  wire pp_4_26_1;
  wire pp_4_27_0;
  wire pp_4_27_1;
  wire pp_4_28_0;
  wire pp_4_28_1;
  wire pp_4_29_0;
  wire pp_4_29_1;
  wire pp_4_30_0;
  wire pp_4_30_1;
  wire pp_4_31_0;
  wire pp_4_31_1;
  assign pp_0_0_0 = pp_0_0;
  assign pp_0_0_1 = be_c_0;
  assign pp_0_1_0 = pp_0_1;
  assign pp_0_2_0 = pp_0_2;
  assign pp_0_2_1 = pp_1_2;
  assign pp_0_2_2 = be_c_1;
  assign pp_0_3_0 = pp_0_3;
  assign pp_0_3_1 = pp_1_3;
  assign pp_0_4_0 = pp_0_4;
  assign pp_0_4_1 = pp_1_4;
  assign pp_0_4_2 = pp_2_4;
  assign pp_0_4_3 = be_c_2;
  assign pp_0_5_0 = pp_0_5;
  assign pp_0_5_1 = pp_1_5;
  assign pp_0_5_2 = pp_2_5;
  assign pp_0_6_0 = pp_0_6;
  assign pp_0_6_1 = pp_1_6;
  assign pp_0_6_2 = pp_2_6;
  assign pp_0_6_3 = pp_3_6;
  assign pp_0_6_4 = be_c_3;
  assign pp_0_7_0 = pp_0_7;
  assign pp_0_7_1 = pp_1_7;
  assign pp_0_7_2 = pp_2_7;
  assign pp_0_7_3 = pp_3_7;
  assign pp_0_8_0 = pp_0_8;
  assign pp_0_8_1 = pp_1_8;
  assign pp_0_8_2 = pp_2_8;
  assign pp_0_8_3 = pp_3_8;
  assign pp_0_8_4 = pp_4_8;
  assign pp_0_8_5 = be_c_4;
  assign pp_0_9_0 = pp_0_9;
  assign pp_0_9_1 = pp_1_9;
  assign pp_0_9_2 = pp_2_9;
  assign pp_0_9_3 = pp_3_9;
  assign pp_0_9_4 = pp_4_9;
  assign pp_0_10_0 = pp_0_10;
  assign pp_0_10_1 = pp_1_10;
  assign pp_0_10_2 = pp_2_10;
  assign pp_0_10_3 = pp_3_10;
  assign pp_0_10_4 = pp_4_10;
  assign pp_0_10_5 = pp_5_10;
  assign pp_0_10_6 = be_c_5;
  assign pp_0_11_0 = pp_0_11;
  assign pp_0_11_1 = pp_1_11;
  assign pp_0_11_2 = pp_2_11;
  assign pp_0_11_3 = pp_3_11;
  assign pp_0_11_4 = pp_4_11;
  assign pp_0_11_5 = pp_5_11;
  assign pp_0_12_0 = pp_0_12;
  assign pp_0_12_1 = pp_1_12;
  assign pp_0_12_2 = pp_2_12;
  assign pp_0_12_3 = pp_3_12;
  assign pp_0_12_4 = pp_4_12;
  assign pp_0_12_5 = pp_5_12;
  assign pp_0_12_6 = pp_6_12;
  assign pp_0_12_7 = be_c_6;
  assign pp_0_13_0 = pp_0_13;
  assign pp_0_13_1 = pp_1_13;
  assign pp_0_13_2 = pp_2_13;
  assign pp_0_13_3 = pp_3_13;
  assign pp_0_13_4 = pp_4_13;
  assign pp_0_13_5 = pp_5_13;
  assign pp_0_13_6 = pp_6_13;
  assign pp_0_14_0 = pp_0_14;
  assign pp_0_14_1 = pp_1_14;
  assign pp_0_14_2 = pp_2_14;
  assign pp_0_14_3 = pp_3_14;
  assign pp_0_14_4 = pp_4_14;
  assign pp_0_14_5 = pp_5_14;
  assign pp_0_14_6 = pp_6_14;
  assign pp_0_14_7 = pp_7_14;
  assign pp_0_14_8 = be_c_7;
  assign pp_0_15_0 = pp_0_15;
  assign pp_0_15_1 = pp_1_15;
  assign pp_0_15_2 = pp_2_15;
  assign pp_0_15_3 = pp_3_15;
  assign pp_0_15_4 = pp_4_15;
  assign pp_0_15_5 = pp_5_15;
  assign pp_0_15_6 = pp_6_15;
  assign pp_0_15_7 = pp_7_15;
  assign pp_0_16_0 = pp_0_16;
  assign pp_0_16_1 = pp_1_16;
  assign pp_0_16_2 = pp_2_16;
  assign pp_0_16_3 = pp_3_16;
  assign pp_0_16_4 = pp_4_16;
  assign pp_0_16_5 = pp_5_16;
  assign pp_0_16_6 = pp_6_16;
  assign pp_0_16_7 = pp_7_16;
  assign pp_0_16_8 = pp_8_16;
  assign pp_0_17_0 = pp_0_17;
  assign pp_0_17_1 = pp_1_17;
  assign pp_0_17_2 = pp_2_17;
  assign pp_0_17_3 = pp_3_17;
  assign pp_0_17_4 = pp_4_17;
  assign pp_0_17_5 = pp_5_17;
  assign pp_0_17_6 = pp_6_17;
  assign pp_0_17_7 = pp_7_17;
  assign pp_0_17_8 = pp_8_17;
  assign pp_0_18_0 = pp_0_17;
  assign pp_0_18_1 = pp_1_18;
  assign pp_0_18_2 = pp_2_18;
  assign pp_0_18_3 = pp_3_18;
  assign pp_0_18_4 = pp_4_18;
  assign pp_0_18_5 = pp_5_18;
  assign pp_0_18_6 = pp_6_18;
  assign pp_0_18_7 = pp_7_18;
  assign pp_0_18_8 = pp_8_18;
  assign pp_0_19_0 = not_pp_0_19;
  assign pp_0_19_1 = not_pp_1_19;
  assign pp_0_19_2 = pp_2_19;
  assign pp_0_19_3 = pp_3_19;
  assign pp_0_19_4 = pp_4_19;
  assign pp_0_19_5 = pp_5_19;
  assign pp_0_19_6 = pp_6_19;
  assign pp_0_19_7 = pp_7_19;
  assign pp_0_19_8 = pp_8_19;
  assign pp_0_20_0 = one;
  assign pp_0_20_1 = pp_2_20;
  assign pp_0_20_2 = pp_3_20;
  assign pp_0_20_3 = pp_4_20;
  assign pp_0_20_4 = pp_5_20;
  assign pp_0_20_5 = pp_6_20;
  assign pp_0_20_6 = pp_7_20;
  assign pp_0_20_7 = pp_8_20;
  assign pp_0_21_0 = not_pp_2_21;
  assign pp_0_21_1 = pp_3_21;
  assign pp_0_21_2 = pp_4_21;
  assign pp_0_21_3 = pp_5_21;
  assign pp_0_21_4 = pp_6_21;
  assign pp_0_21_5 = pp_7_21;
  assign pp_0_21_6 = pp_8_21;
  assign pp_0_22_0 = one;
  assign pp_0_22_1 = pp_3_22;
  assign pp_0_22_2 = pp_4_22;
  assign pp_0_22_3 = pp_5_22;
  assign pp_0_22_4 = pp_6_22;
  assign pp_0_22_5 = pp_7_22;
  assign pp_0_22_6 = pp_8_22;
  assign pp_0_23_0 = not_pp_3_23;
  assign pp_0_23_1 = pp_4_23;
  assign pp_0_23_2 = pp_5_23;
  assign pp_0_23_3 = pp_6_23;
  assign pp_0_23_4 = pp_7_23;
  assign pp_0_23_5 = pp_8_23;
  assign pp_0_24_0 = one;
  assign pp_0_24_1 = pp_4_24;
  assign pp_0_24_2 = pp_5_24;
  assign pp_0_24_3 = pp_6_24;
  assign pp_0_24_4 = pp_7_24;
  assign pp_0_24_5 = pp_8_24;
  assign pp_0_25_0 = not_pp_4_25;
  assign pp_0_25_1 = pp_5_25;
  assign pp_0_25_2 = pp_6_25;
  assign pp_0_25_3 = pp_7_25;
  assign pp_0_25_4 = pp_8_25;
  assign pp_0_26_0 = one;
  assign pp_0_26_1 = pp_5_26;
  assign pp_0_26_2 = pp_6_26;
  assign pp_0_26_3 = pp_7_26;
  assign pp_0_26_4 = pp_8_26;
  assign pp_0_27_0 = not_pp_5_27;
  assign pp_0_27_1 = pp_6_27;
  assign pp_0_27_2 = pp_7_27;
  assign pp_0_27_3 = pp_8_27;
  assign pp_0_28_0 = one;
  assign pp_0_28_1 = pp_6_28;
  assign pp_0_28_2 = pp_7_28;
  assign pp_0_28_3 = pp_8_28;
  assign pp_0_29_0 = not_pp_6_29;
  assign pp_0_29_1 = pp_7_29;
  assign pp_0_29_2 = pp_8_29;
  assign pp_0_30_0 = one;
  assign pp_0_30_1 = pp_7_30;
  assign pp_0_30_2 = pp_8_30;
  assign pp_0_31_0 = not_pp_7_31;
  assign pp_0_31_1 = pp_8_31;

  assign pp_1_0_0 = pp_0_0_0;
  assign pp_1_0_1 = pp_0_0_1;
  assign pp_1_1_0 = pp_0_1_0;
  assign pp_1_2_0 = pp_0_2_0;
  assign pp_1_2_1 = pp_0_2_1;
  assign pp_1_2_2 = pp_0_2_2;
  MG_HA ha_0_3_0(
    .a(pp_0_3_0),
    .b(pp_0_3_1),
    .sum(pp_1_3_0),
    .cout(pp_1_4_0)
  );

  assign pp_1_4_1 = pp_0_4_0;
  assign pp_1_4_2 = pp_0_4_1;
  assign pp_1_4_3 = pp_0_4_2;
  assign pp_1_4_4 = pp_0_4_3;
  MG_FA fa_0_5_0(
    .a(pp_0_5_0),
    .b(pp_0_5_1),
    .cin(pp_0_5_2),
    .sum(pp_1_5_0),
    .cout(pp_1_6_0)
  );

  MG_FA fa_0_6_0(
    .a(pp_0_6_0),
    .b(pp_0_6_1),
    .cin(pp_0_6_2),
    .sum(pp_1_6_1),
    .cout(pp_1_7_0)
  );

  MG_HA ha_0_6_1(
    .a(pp_0_6_3),
    .b(pp_0_6_4),
    .sum(pp_1_6_2),
    .cout(pp_1_7_1)
  );

  MG_FA fa_0_7_0(
    .a(pp_0_7_0),
    .b(pp_0_7_1),
    .cin(pp_0_7_2),
    .sum(pp_1_7_2),
    .cout(pp_1_8_0)
  );

  assign pp_1_7_3 = pp_0_7_3;
  MG_FA fa_0_8_0(
    .a(pp_0_8_0),
    .b(pp_0_8_1),
    .cin(pp_0_8_2),
    .sum(pp_1_8_1),
    .cout(pp_1_9_0)
  );

  MG_FA fa_0_8_1(
    .a(pp_0_8_3),
    .b(pp_0_8_4),
    .cin(pp_0_8_5),
    .sum(pp_1_8_2),
    .cout(pp_1_9_1)
  );

  MG_FA fa_0_9_0(
    .a(pp_0_9_0),
    .b(pp_0_9_1),
    .cin(pp_0_9_2),
    .sum(pp_1_9_2),
    .cout(pp_1_10_0)
  );

  assign pp_1_9_3 = pp_0_9_3;
  assign pp_1_9_4 = pp_0_9_4;
  MG_FA fa_0_10_0(
    .a(pp_0_10_0),
    .b(pp_0_10_1),
    .cin(pp_0_10_2),
    .sum(pp_1_10_1),
    .cout(pp_1_11_0)
  );

  MG_FA fa_0_10_1(
    .a(pp_0_10_3),
    .b(pp_0_10_4),
    .cin(pp_0_10_5),
    .sum(pp_1_10_2),
    .cout(pp_1_11_1)
  );

  assign pp_1_10_3 = pp_0_10_6;
  MG_FA fa_0_11_0(
    .a(pp_0_11_0),
    .b(pp_0_11_1),
    .cin(pp_0_11_2),
    .sum(pp_1_11_2),
    .cout(pp_1_12_0)
  );

  assign pp_1_11_3 = pp_0_11_3;
  assign pp_1_11_4 = pp_0_11_4;
  assign pp_1_11_5 = pp_0_11_5;
  MG_FA fa_0_12_0(
    .a(pp_0_12_0),
    .b(pp_0_12_1),
    .cin(pp_0_12_2),
    .sum(pp_1_12_1),
    .cout(pp_1_13_0)
  );

  MG_FA fa_0_12_1(
    .a(pp_0_12_3),
    .b(pp_0_12_4),
    .cin(pp_0_12_5),
    .sum(pp_1_12_2),
    .cout(pp_1_13_1)
  );

  MG_HA ha_0_12_2(
    .a(pp_0_12_6),
    .b(pp_0_12_7),
    .sum(pp_1_12_3),
    .cout(pp_1_13_2)
  );

  MG_FA fa_0_13_0(
    .a(pp_0_13_0),
    .b(pp_0_13_1),
    .cin(pp_0_13_2),
    .sum(pp_1_13_3),
    .cout(pp_1_14_0)
  );

  MG_FA fa_0_13_1(
    .a(pp_0_13_3),
    .b(pp_0_13_4),
    .cin(pp_0_13_5),
    .sum(pp_1_13_4),
    .cout(pp_1_14_1)
  );

  assign pp_1_13_5 = pp_0_13_6;
  MG_FA fa_0_14_0(
    .a(pp_0_14_0),
    .b(pp_0_14_1),
    .cin(pp_0_14_2),
    .sum(pp_1_14_2),
    .cout(pp_1_15_0)
  );

  MG_FA fa_0_14_1(
    .a(pp_0_14_3),
    .b(pp_0_14_4),
    .cin(pp_0_14_5),
    .sum(pp_1_14_3),
    .cout(pp_1_15_1)
  );

  MG_HA ha_0_14_2(
    .a(pp_0_14_6),
    .b(pp_0_14_7),
    .sum(pp_1_14_4),
    .cout(pp_1_15_2)
  );

  assign pp_1_14_5 = pp_0_14_8;
  MG_FA fa_0_15_0(
    .a(pp_0_15_0),
    .b(pp_0_15_1),
    .cin(pp_0_15_2),
    .sum(pp_1_15_3),
    .cout(pp_1_16_0)
  );

  MG_FA fa_0_15_1(
    .a(pp_0_15_3),
    .b(pp_0_15_4),
    .cin(pp_0_15_5),
    .sum(pp_1_15_4),
    .cout(pp_1_16_1)
  );

  MG_HA ha_0_15_2(
    .a(pp_0_15_6),
    .b(pp_0_15_7),
    .sum(pp_1_15_5),
    .cout(pp_1_16_2)
  );

  MG_FA fa_0_16_0(
    .a(pp_0_16_0),
    .b(pp_0_16_1),
    .cin(pp_0_16_2),
    .sum(pp_1_16_3),
    .cout(pp_1_17_0)
  );

  MG_FA fa_0_16_1(
    .a(pp_0_16_3),
    .b(pp_0_16_4),
    .cin(pp_0_16_5),
    .sum(pp_1_16_4),
    .cout(pp_1_17_1)
  );

  MG_FA fa_0_16_2(
    .a(pp_0_16_6),
    .b(pp_0_16_7),
    .cin(pp_0_16_8),
    .sum(pp_1_16_5),
    .cout(pp_1_17_2)
  );

  MG_FA fa_0_17_0(
    .a(pp_0_17_0),
    .b(pp_0_17_1),
    .cin(pp_0_17_2),
    .sum(pp_1_17_3),
    .cout(pp_1_18_0)
  );

  MG_FA fa_0_17_1(
    .a(pp_0_17_3),
    .b(pp_0_17_4),
    .cin(pp_0_17_5),
    .sum(pp_1_17_4),
    .cout(pp_1_18_1)
  );

  MG_FA fa_0_17_2(
    .a(pp_0_17_6),
    .b(pp_0_17_7),
    .cin(pp_0_17_8),
    .sum(pp_1_17_5),
    .cout(pp_1_18_2)
  );

  MG_FA fa_0_18_0(
    .a(pp_0_18_0),
    .b(pp_0_18_1),
    .cin(pp_0_18_2),
    .sum(pp_1_18_3),
    .cout(pp_1_19_0)
  );

  MG_FA fa_0_18_1(
    .a(pp_0_18_3),
    .b(pp_0_18_4),
    .cin(pp_0_18_5),
    .sum(pp_1_18_4),
    .cout(pp_1_19_1)
  );

  MG_FA fa_0_18_2(
    .a(pp_0_18_6),
    .b(pp_0_18_7),
    .cin(pp_0_18_8),
    .sum(pp_1_18_5),
    .cout(pp_1_19_2)
  );

  MG_FA fa_0_19_0(
    .a(pp_0_19_0),
    .b(pp_0_19_1),
    .cin(pp_0_19_2),
    .sum(pp_1_19_3),
    .cout(pp_1_20_0)
  );

  MG_FA fa_0_19_1(
    .a(pp_0_19_3),
    .b(pp_0_19_4),
    .cin(pp_0_19_5),
    .sum(pp_1_19_4),
    .cout(pp_1_20_1)
  );

  MG_FA fa_0_19_2(
    .a(pp_0_19_6),
    .b(pp_0_19_7),
    .cin(pp_0_19_8),
    .sum(pp_1_19_5),
    .cout(pp_1_20_2)
  );

  MG_FA fa_0_20_0(
    .a(pp_0_20_0),
    .b(pp_0_20_1),
    .cin(pp_0_20_2),
    .sum(pp_1_20_3),
    .cout(pp_1_21_0)
  );

  MG_FA fa_0_20_1(
    .a(pp_0_20_3),
    .b(pp_0_20_4),
    .cin(pp_0_20_5),
    .sum(pp_1_20_4),
    .cout(pp_1_21_1)
  );

  MG_HA ha_0_20_2(
    .a(pp_0_20_6),
    .b(pp_0_20_7),
    .sum(pp_1_20_5),
    .cout(pp_1_21_2)
  );

  MG_FA fa_0_21_0(
    .a(pp_0_21_0),
    .b(pp_0_21_1),
    .cin(pp_0_21_2),
    .sum(pp_1_21_3),
    .cout(pp_1_22_0)
  );

  MG_FA fa_0_21_1(
    .a(pp_0_21_3),
    .b(pp_0_21_4),
    .cin(pp_0_21_5),
    .sum(pp_1_21_4),
    .cout(pp_1_22_1)
  );

  assign pp_1_21_5 = pp_0_21_6;
  MG_FA fa_0_22_0(
    .a(pp_0_22_0),
    .b(pp_0_22_1),
    .cin(pp_0_22_2),
    .sum(pp_1_22_2),
    .cout(pp_1_23_0)
  );

  MG_HA ha_0_22_1(
    .a(pp_0_22_3),
    .b(pp_0_22_4),
    .sum(pp_1_22_3),
    .cout(pp_1_23_1)
  );

  assign pp_1_22_4 = pp_0_22_5;
  assign pp_1_22_5 = pp_0_22_6;
  MG_FA fa_0_23_0(
    .a(pp_0_23_0),
    .b(pp_0_23_1),
    .cin(pp_0_23_2),
    .sum(pp_1_23_2),
    .cout(pp_1_24_0)
  );

  MG_FA fa_0_23_1(
    .a(pp_0_23_3),
    .b(pp_0_23_4),
    .cin(pp_0_23_5),
    .sum(pp_1_23_3),
    .cout(pp_1_24_1)
  );

  MG_FA fa_0_24_0(
    .a(pp_0_24_0),
    .b(pp_0_24_1),
    .cin(pp_0_24_2),
    .sum(pp_1_24_2),
    .cout(pp_1_25_0)
  );

  assign pp_1_24_3 = pp_0_24_3;
  assign pp_1_24_4 = pp_0_24_4;
  assign pp_1_24_5 = pp_0_24_5;
  assign pp_1_25_1 = pp_0_25_0;
  assign pp_1_25_2 = pp_0_25_1;
  assign pp_1_25_3 = pp_0_25_2;
  assign pp_1_25_4 = pp_0_25_3;
  assign pp_1_25_5 = pp_0_25_4;
  MG_FA fa_0_26_0(
    .a(pp_0_26_0),
    .b(pp_0_26_1),
    .cin(pp_0_26_2),
    .sum(pp_1_26_0),
    .cout(pp_1_27_0)
  );

  assign pp_1_26_1 = pp_0_26_3;
  assign pp_1_26_2 = pp_0_26_4;
  MG_FA fa_0_27_0(
    .a(pp_0_27_0),
    .b(pp_0_27_1),
    .cin(pp_0_27_2),
    .sum(pp_1_27_1),
    .cout(pp_1_28_0)
  );

  assign pp_1_27_2 = pp_0_27_3;
  MG_FA fa_0_28_0(
    .a(pp_0_28_0),
    .b(pp_0_28_1),
    .cin(pp_0_28_2),
    .sum(pp_1_28_1),
    .cout(pp_1_29_0)
  );

  assign pp_1_28_2 = pp_0_28_3;
  assign pp_1_29_1 = pp_0_29_0;
  assign pp_1_29_2 = pp_0_29_1;
  assign pp_1_29_3 = pp_0_29_2;
  assign pp_1_30_0 = pp_0_30_0;
  assign pp_1_30_1 = pp_0_30_1;
  assign pp_1_30_2 = pp_0_30_2;
  assign pp_1_31_0 = pp_0_31_0;
  assign pp_1_31_1 = pp_0_31_1;
  assign pp_2_0_0 = pp_1_0_0;
  assign pp_2_0_1 = pp_1_0_1;
  assign pp_2_1_0 = pp_1_1_0;
  assign pp_2_2_0 = pp_1_2_0;
  assign pp_2_2_1 = pp_1_2_1;
  assign pp_2_2_2 = pp_1_2_2;
  assign pp_2_3_0 = pp_1_3_0;
  MG_FA fa_1_4_0(
    .a(pp_1_4_0),
    .b(pp_1_4_1),
    .cin(pp_1_4_2),
    .sum(pp_2_4_0),
    .cout(pp_2_5_0)
  );

  assign pp_2_4_1 = pp_1_4_3;
  assign pp_2_4_2 = pp_1_4_4;
  assign pp_2_5_1 = pp_1_5_0;
  MG_FA fa_1_6_0(
    .a(pp_1_6_0),
    .b(pp_1_6_1),
    .cin(pp_1_6_2),
    .sum(pp_2_6_0),
    .cout(pp_2_7_0)
  );

  MG_FA fa_1_7_0(
    .a(pp_1_7_0),
    .b(pp_1_7_1),
    .cin(pp_1_7_2),
    .sum(pp_2_7_1),
    .cout(pp_2_8_0)
  );

  assign pp_2_7_2 = pp_1_7_3;
  MG_FA fa_1_8_0(
    .a(pp_1_8_0),
    .b(pp_1_8_1),
    .cin(pp_1_8_2),
    .sum(pp_2_8_1),
    .cout(pp_2_9_0)
  );

  MG_FA fa_1_9_0(
    .a(pp_1_9_0),
    .b(pp_1_9_1),
    .cin(pp_1_9_2),
    .sum(pp_2_9_1),
    .cout(pp_2_10_0)
  );

  assign pp_2_9_2 = pp_1_9_3;
  assign pp_2_9_3 = pp_1_9_4;
  MG_FA fa_1_10_0(
    .a(pp_1_10_0),
    .b(pp_1_10_1),
    .cin(pp_1_10_2),
    .sum(pp_2_10_1),
    .cout(pp_2_11_0)
  );

  assign pp_2_10_2 = pp_1_10_3;
  MG_FA fa_1_11_0(
    .a(pp_1_11_0),
    .b(pp_1_11_1),
    .cin(pp_1_11_2),
    .sum(pp_2_11_1),
    .cout(pp_2_12_0)
  );

  MG_FA fa_1_11_1(
    .a(pp_1_11_3),
    .b(pp_1_11_4),
    .cin(pp_1_11_5),
    .sum(pp_2_11_2),
    .cout(pp_2_12_1)
  );

  assign pp_2_12_2 = pp_1_12_0;
  assign pp_2_12_3 = pp_1_12_1;
  assign pp_2_12_4 = pp_1_12_2;
  assign pp_2_12_5 = pp_1_12_3;
  MG_FA fa_1_13_0(
    .a(pp_1_13_0),
    .b(pp_1_13_1),
    .cin(pp_1_13_2),
    .sum(pp_2_13_0),
    .cout(pp_2_14_0)
  );

  MG_FA fa_1_13_1(
    .a(pp_1_13_3),
    .b(pp_1_13_4),
    .cin(pp_1_13_5),
    .sum(pp_2_13_1),
    .cout(pp_2_14_1)
  );

  MG_FA fa_1_14_0(
    .a(pp_1_14_0),
    .b(pp_1_14_1),
    .cin(pp_1_14_2),
    .sum(pp_2_14_2),
    .cout(pp_2_15_0)
  );

  MG_FA fa_1_14_1(
    .a(pp_1_14_3),
    .b(pp_1_14_4),
    .cin(pp_1_14_5),
    .sum(pp_2_14_3),
    .cout(pp_2_15_1)
  );

  MG_FA fa_1_15_0(
    .a(pp_1_15_0),
    .b(pp_1_15_1),
    .cin(pp_1_15_2),
    .sum(pp_2_15_2),
    .cout(pp_2_16_0)
  );

  assign pp_2_15_3 = pp_1_15_3;
  assign pp_2_15_4 = pp_1_15_4;
  assign pp_2_15_5 = pp_1_15_5;
  MG_FA fa_1_16_0(
    .a(pp_1_16_0),
    .b(pp_1_16_1),
    .cin(pp_1_16_2),
    .sum(pp_2_16_1),
    .cout(pp_2_17_0)
  );

  MG_FA fa_1_16_1(
    .a(pp_1_16_3),
    .b(pp_1_16_4),
    .cin(pp_1_16_5),
    .sum(pp_2_16_2),
    .cout(pp_2_17_1)
  );

  MG_FA fa_1_17_0(
    .a(pp_1_17_0),
    .b(pp_1_17_1),
    .cin(pp_1_17_2),
    .sum(pp_2_17_2),
    .cout(pp_2_18_0)
  );

  MG_FA fa_1_17_1(
    .a(pp_1_17_3),
    .b(pp_1_17_4),
    .cin(pp_1_17_5),
    .sum(pp_2_17_3),
    .cout(pp_2_18_1)
  );

  MG_FA fa_1_18_0(
    .a(pp_1_18_0),
    .b(pp_1_18_1),
    .cin(pp_1_18_2),
    .sum(pp_2_18_2),
    .cout(pp_2_19_0)
  );

  assign pp_2_18_3 = pp_1_18_3;
  assign pp_2_18_4 = pp_1_18_4;
  assign pp_2_18_5 = pp_1_18_5;
  MG_FA fa_1_19_0(
    .a(pp_1_19_0),
    .b(pp_1_19_1),
    .cin(pp_1_19_2),
    .sum(pp_2_19_1),
    .cout(pp_2_20_0)
  );

  MG_FA fa_1_19_1(
    .a(pp_1_19_3),
    .b(pp_1_19_4),
    .cin(pp_1_19_5),
    .sum(pp_2_19_2),
    .cout(pp_2_20_1)
  );

  MG_FA fa_1_20_0(
    .a(pp_1_20_0),
    .b(pp_1_20_1),
    .cin(pp_1_20_2),
    .sum(pp_2_20_2),
    .cout(pp_2_21_0)
  );

  MG_FA fa_1_20_1(
    .a(pp_1_20_3),
    .b(pp_1_20_4),
    .cin(pp_1_20_5),
    .sum(pp_2_20_3),
    .cout(pp_2_21_1)
  );

  MG_FA fa_1_21_0(
    .a(pp_1_21_0),
    .b(pp_1_21_1),
    .cin(pp_1_21_2),
    .sum(pp_2_21_2),
    .cout(pp_2_22_0)
  );

  MG_FA fa_1_21_1(
    .a(pp_1_21_3),
    .b(pp_1_21_4),
    .cin(pp_1_21_5),
    .sum(pp_2_21_3),
    .cout(pp_2_22_1)
  );

  MG_FA fa_1_22_0(
    .a(pp_1_22_0),
    .b(pp_1_22_1),
    .cin(pp_1_22_2),
    .sum(pp_2_22_2),
    .cout(pp_2_23_0)
  );

  MG_FA fa_1_22_1(
    .a(pp_1_22_3),
    .b(pp_1_22_4),
    .cin(pp_1_22_5),
    .sum(pp_2_22_3),
    .cout(pp_2_23_1)
  );

  MG_FA fa_1_23_0(
    .a(pp_1_23_0),
    .b(pp_1_23_1),
    .cin(pp_1_23_2),
    .sum(pp_2_23_2),
    .cout(pp_2_24_0)
  );

  assign pp_2_23_3 = pp_1_23_3;
  MG_HA ha_1_24_0(
    .a(pp_1_24_0),
    .b(pp_1_24_1),
    .sum(pp_2_24_1),
    .cout(pp_2_25_0)
  );

  assign pp_2_24_2 = pp_1_24_2;
  assign pp_2_24_3 = pp_1_24_3;
  assign pp_2_24_4 = pp_1_24_4;
  assign pp_2_24_5 = pp_1_24_5;
  MG_FA fa_1_25_0(
    .a(pp_1_25_0),
    .b(pp_1_25_1),
    .cin(pp_1_25_2),
    .sum(pp_2_25_1),
    .cout(pp_2_26_0)
  );

  MG_FA fa_1_25_1(
    .a(pp_1_25_3),
    .b(pp_1_25_4),
    .cin(pp_1_25_5),
    .sum(pp_2_25_2),
    .cout(pp_2_26_1)
  );

  MG_FA fa_1_26_0(
    .a(pp_1_26_0),
    .b(pp_1_26_1),
    .cin(pp_1_26_2),
    .sum(pp_2_26_2),
    .cout(pp_2_27_0)
  );

  MG_FA fa_1_27_0(
    .a(pp_1_27_0),
    .b(pp_1_27_1),
    .cin(pp_1_27_2),
    .sum(pp_2_27_1),
    .cout(pp_2_28_0)
  );

  MG_FA fa_1_28_0(
    .a(pp_1_28_0),
    .b(pp_1_28_1),
    .cin(pp_1_28_2),
    .sum(pp_2_28_1),
    .cout(pp_2_29_0)
  );

  MG_FA fa_1_29_0(
    .a(pp_1_29_0),
    .b(pp_1_29_1),
    .cin(pp_1_29_2),
    .sum(pp_2_29_1),
    .cout(pp_2_30_0)
  );

  assign pp_2_29_2 = pp_1_29_3;
  MG_FA fa_1_30_0(
    .a(pp_1_30_0),
    .b(pp_1_30_1),
    .cin(pp_1_30_2),
    .sum(pp_2_30_1),
    .cout(pp_2_31_0)
  );

  assign pp_2_31_1 = pp_1_31_0;
  assign pp_2_31_2 = pp_1_31_1;
  assign pp_3_0_0 = pp_2_0_0;
  assign pp_3_0_1 = pp_2_0_1;
  assign pp_3_1_0 = pp_2_1_0;
  MG_HA ha_2_2_0(
    .a(pp_2_2_0),
    .b(pp_2_2_1),
    .sum(pp_3_2_0),
    .cout(pp_3_3_0)
  );

  assign pp_3_2_1 = pp_2_2_2;
  assign pp_3_3_1 = pp_2_3_0;
  MG_HA ha_2_4_0(
    .a(pp_2_4_0),
    .b(pp_2_4_1),
    .sum(pp_3_4_0),
    .cout(pp_3_5_0)
  );

  assign pp_3_4_1 = pp_2_4_2;
  assign pp_3_5_1 = pp_2_5_0;
  assign pp_3_5_2 = pp_2_5_1;
  assign pp_3_6_0 = pp_2_6_0;
  MG_HA ha_2_7_0(
    .a(pp_2_7_0),
    .b(pp_2_7_1),
    .sum(pp_3_7_0),
    .cout(pp_3_8_0)
  );

  assign pp_3_7_1 = pp_2_7_2;
  MG_HA ha_2_8_0(
    .a(pp_2_8_0),
    .b(pp_2_8_1),
    .sum(pp_3_8_1),
    .cout(pp_3_9_0)
  );

  MG_FA fa_2_9_0(
    .a(pp_2_9_0),
    .b(pp_2_9_1),
    .cin(pp_2_9_2),
    .sum(pp_3_9_1),
    .cout(pp_3_10_0)
  );

  assign pp_3_9_2 = pp_2_9_3;
  MG_HA ha_2_10_0(
    .a(pp_2_10_0),
    .b(pp_2_10_2),
    .sum(pp_3_10_1),
    .cout(pp_3_11_0)
  );

  assign pp_3_10_2 = pp_2_10_1;
  MG_HA ha_2_11_0(
    .a(pp_2_11_0),
    .b(pp_2_11_1),
    .sum(pp_3_11_1),
    .cout(pp_3_12_0)
  );

  assign pp_3_11_2 = pp_2_11_2;
  MG_FA fa_2_12_0(
    .a(pp_2_12_2),
    .b(pp_2_12_1),
    .cin(pp_2_12_0),
    .sum(pp_3_12_1),
    .cout(pp_3_13_0)
  );

  MG_FA fa_2_12_1(
    .a(pp_2_12_3),
    .b(pp_2_12_4),
    .cin(pp_2_12_5),
    .sum(pp_3_12_2),
    .cout(pp_3_13_1)
  );

  MG_HA ha_2_13_0(
    .a(pp_2_13_0),
    .b(pp_2_13_1),
    .sum(pp_3_13_2),
    .cout(pp_3_14_0)
  );

  MG_FA fa_2_14_0(
    .a(pp_2_14_0),
    .b(pp_2_14_1),
    .cin(pp_2_14_2),
    .sum(pp_3_14_1),
    .cout(pp_3_15_0)
  );

  assign pp_3_14_2 = pp_2_14_3;
  MG_FA fa_2_15_0(
    .a(pp_2_15_5),
    .b(pp_2_15_1),
    .cin(pp_2_15_2),
    .sum(pp_3_15_1),
    .cout(pp_3_16_0)
  );

  MG_FA fa_2_15_1(
    .a(pp_2_15_3),
    .b(pp_2_15_4),
    .cin(pp_2_15_0),
    .sum(pp_3_15_2),
    .cout(pp_3_16_1)
  );

  MG_FA fa_2_16_0(
    .a(pp_2_16_0),
    .b(pp_2_16_1),
    .cin(pp_2_16_2),
    .sum(pp_3_16_2),
    .cout(pp_3_17_0)
  );

  MG_FA fa_2_17_0(
    .a(pp_2_17_0),
    .b(pp_2_17_1),
    .cin(pp_2_17_2),
    .sum(pp_3_17_1),
    .cout(pp_3_18_0)
  );

  assign pp_3_17_2 = pp_2_17_3;
  MG_FA fa_2_18_0(
    .a(pp_2_18_0),
    .b(pp_2_18_1),
    .cin(pp_2_18_2),
    .sum(pp_3_18_1),
    .cout(pp_3_19_0)
  );

  MG_FA fa_2_18_1(
    .a(pp_2_18_3),
    .b(pp_2_18_4),
    .cin(pp_2_18_5),
    .sum(pp_3_18_2),
    .cout(pp_3_19_1)
  );

  MG_FA fa_2_19_0(
    .a(pp_2_19_0),
    .b(pp_2_19_1),
    .cin(pp_2_19_2),
    .sum(pp_3_19_2),
    .cout(pp_3_20_0)
  );

  MG_FA fa_2_20_0(
    .a(pp_2_20_0),
    .b(pp_2_20_1),
    .cin(pp_2_20_2),
    .sum(pp_3_20_1),
    .cout(pp_3_21_0)
  );

  assign pp_3_20_2 = pp_2_20_3;
  MG_FA fa_2_21_0(
    .a(pp_2_21_0),
    .b(pp_2_21_1),
    .cin(pp_2_21_2),
    .sum(pp_3_21_1),
    .cout(pp_3_22_0)
  );

  assign pp_3_21_2 = pp_2_21_3;
  MG_FA fa_2_22_0(
    .a(pp_2_22_0),
    .b(pp_2_22_1),
    .cin(pp_2_22_2),
    .sum(pp_3_22_1),
    .cout(pp_3_23_0)
  );

  assign pp_3_22_2 = pp_2_22_3;
  MG_FA fa_2_23_0(
    .a(pp_2_23_3),
    .b(pp_2_23_1),
    .cin(pp_2_23_2),
    .sum(pp_3_23_1),
    .cout(pp_3_24_0)
  );

  assign pp_3_23_2 = pp_2_23_0;
  MG_FA fa_2_24_0(
    .a(pp_2_24_3),
    .b(pp_2_24_1),
    .cin(pp_2_24_2),
    .sum(pp_3_24_1),
    .cout(pp_3_25_0)
  );

  MG_FA fa_2_24_1(
    .a(pp_2_24_0),
    .b(pp_2_24_4),
    .cin(pp_2_24_5),
    .sum(pp_3_24_2),
    .cout(pp_3_25_1)
  );

  MG_FA fa_2_25_0(
    .a(pp_2_25_0),
    .b(pp_2_25_1),
    .cin(pp_2_25_2),
    .sum(pp_3_25_2),
    .cout(pp_3_26_0)
  );

  MG_HA ha_2_26_0(
    .a(pp_2_26_0),
    .b(pp_2_26_1),
    .sum(pp_3_26_1),
    .cout(pp_3_27_0)
  );

  assign pp_3_26_2 = pp_2_26_2;
  assign pp_3_27_1 = pp_2_27_0;
  assign pp_3_27_2 = pp_2_27_1;
  MG_HA ha_2_28_0(
    .a(pp_2_28_0),
    .b(pp_2_28_1),
    .sum(pp_3_28_0),
    .cout(pp_3_29_0)
  );

  MG_FA fa_2_29_0(
    .a(pp_2_29_0),
    .b(pp_2_29_1),
    .cin(pp_2_29_2),
    .sum(pp_3_29_1),
    .cout(pp_3_30_0)
  );

  assign pp_3_30_1 = pp_2_30_0;
  assign pp_3_30_2 = pp_2_30_1;
  MG_FA fa_2_31_0(
    .a(pp_2_31_0),
    .b(pp_2_31_1),
    .cin(pp_2_31_2),
    .sum(pp_3_31_0),
    .cout()
  );

  assign pp_4_0_0 = pp_3_0_0;
  assign pp_4_0_1 = pp_3_0_1;
  assign pp_4_1_0 = pp_3_1_0;
  assign pp_4_2_0 = pp_3_2_0;
  assign pp_4_2_1 = pp_3_2_1;
  assign pp_4_3_0 = pp_3_3_0;
  assign pp_4_3_1 = pp_3_3_1;
  assign pp_4_4_0 = pp_3_4_0;
  assign pp_4_4_1 = pp_3_4_1;
  MG_HA ha_3_5_0(
    .a(pp_3_5_0),
    .b(pp_3_5_1),
    .sum(pp_4_5_0),
    .cout(pp_4_6_0)
  );

  assign pp_4_5_1 = pp_3_5_2;
  assign pp_4_6_1 = pp_3_6_0;
  assign pp_4_7_0 = pp_3_7_0;
  assign pp_4_7_1 = pp_3_7_1;
  assign pp_4_8_0 = pp_3_8_0;
  assign pp_4_8_1 = pp_3_8_1;
  MG_HA ha_3_9_0(
    .a(pp_3_9_0),
    .b(pp_3_9_1),
    .sum(pp_4_9_0),
    .cout(pp_4_10_0)
  );

  assign pp_4_9_1 = pp_3_9_2;
  MG_FA fa_3_10_0(
    .a(pp_3_10_0),
    .b(pp_3_10_2),
    .cin(pp_3_10_1),
    .sum(pp_4_10_1),
    .cout(pp_4_11_0)
  );

  MG_FA fa_3_11_0(
    .a(pp_3_11_0),
    .b(pp_3_11_1),
    .cin(pp_3_11_2),
    .sum(pp_4_11_1),
    .cout(pp_4_12_0)
  );

  MG_FA fa_3_12_0(
    .a(pp_3_12_0),
    .b(pp_3_12_1),
    .cin(pp_3_12_2),
    .sum(pp_4_12_1),
    .cout(pp_4_13_0)
  );

  MG_FA fa_3_13_0(
    .a(pp_3_13_0),
    .b(pp_3_13_1),
    .cin(pp_3_13_2),
    .sum(pp_4_13_1),
    .cout(pp_4_14_0)
  );

  MG_FA fa_3_14_0(
    .a(pp_3_14_0),
    .b(pp_3_14_1),
    .cin(pp_3_14_2),
    .sum(pp_4_14_1),
    .cout(pp_4_15_0)
  );

  MG_FA fa_3_15_0(
    .a(pp_3_15_0),
    .b(pp_3_15_1),
    .cin(pp_3_15_2),
    .sum(pp_4_15_1),
    .cout(pp_4_16_0)
  );

  MG_FA fa_3_16_0(
    .a(pp_3_16_0),
    .b(pp_3_16_1),
    .cin(pp_3_16_2),
    .sum(pp_4_16_1),
    .cout(pp_4_17_0)
  );

  MG_FA fa_3_17_0(
    .a(pp_3_17_0),
    .b(pp_3_17_1),
    .cin(pp_3_17_2),
    .sum(pp_4_17_1),
    .cout(pp_4_18_0)
  );

  MG_FA fa_3_18_0(
    .a(pp_3_18_0),
    .b(pp_3_18_1),
    .cin(pp_3_18_2),
    .sum(pp_4_18_1),
    .cout(pp_4_19_0)
  );

  MG_FA fa_3_19_0(
    .a(pp_3_19_0),
    .b(pp_3_19_1),
    .cin(pp_3_19_2),
    .sum(pp_4_19_1),
    .cout(pp_4_20_0)
  );

  MG_FA fa_3_20_0(
    .a(pp_3_20_0),
    .b(pp_3_20_1),
    .cin(pp_3_20_2),
    .sum(pp_4_20_1),
    .cout(pp_4_21_0)
  );

  MG_FA fa_3_21_0(
    .a(pp_3_21_0),
    .b(pp_3_21_1),
    .cin(pp_3_21_2),
    .sum(pp_4_21_1),
    .cout(pp_4_22_0)
  );

  MG_FA fa_3_22_0(
    .a(pp_3_22_0),
    .b(pp_3_22_2),
    .cin(pp_3_22_1),
    .sum(pp_4_22_1),
    .cout(pp_4_23_0)
  );

  MG_FA fa_3_23_0(
    .a(pp_3_23_0),
    .b(pp_3_23_1),
    .cin(pp_3_23_2),
    .sum(pp_4_23_1),
    .cout(pp_4_24_0)
  );

  MG_FA fa_3_24_0(
    .a(pp_3_24_0),
    .b(pp_3_24_1),
    .cin(pp_3_24_2),
    .sum(pp_4_24_1),
    .cout(pp_4_25_0)
  );

  MG_FA fa_3_25_0(
    .a(pp_3_25_0),
    .b(pp_3_25_1),
    .cin(pp_3_25_2),
    .sum(pp_4_25_1),
    .cout(pp_4_26_0)
  );

  MG_FA fa_3_26_0(
    .a(pp_3_26_0),
    .b(pp_3_26_1),
    .cin(pp_3_26_2),
    .sum(pp_4_26_1),
    .cout(pp_4_27_0)
  );

  MG_FA fa_3_27_0(
    .a(pp_3_27_0),
    .b(pp_3_27_1),
    .cin(pp_3_27_2),
    .sum(pp_4_27_1),
    .cout(pp_4_28_0)
  );

  assign pp_4_28_1 = pp_3_28_0;
  assign pp_4_29_0 = pp_3_29_0;
  assign pp_4_29_1 = pp_3_29_1;
  MG_HA ha_3_30_0(
    .a(pp_3_30_0),
    .b(pp_3_30_1),
    .sum(pp_4_30_0),
    .cout(pp_4_31_0)
  );

  assign pp_4_30_1 = pp_3_30_2;
  assign pp_4_31_1 = pp_3_31_0;
  wire [31:0] cta;
  wire [31:0] ctb;
  wire [31:0] cts;
  wire ctc;

  MG_CPA cpa(
 .a(cta), .b(ctb), .sum(cts), .cout(ctc)
  );

  assign cta[0] = pp_4_0_0;
  assign ctb[0] = pp_4_0_1;
  assign cta[1] = pp_4_1_0;
  assign ctb[1] = 1'b0;
  assign cta[2] = pp_4_2_0;
  assign ctb[2] = pp_4_2_1;
  assign cta[3] = pp_4_3_0;
  assign ctb[3] = pp_4_3_1;
  assign cta[4] = pp_4_4_0;
  assign ctb[4] = pp_4_4_1;
  assign cta[5] = pp_4_5_0;
  assign ctb[5] = pp_4_5_1;
  assign cta[6] = pp_4_6_0;
  assign ctb[6] = pp_4_6_1;
  assign cta[7] = pp_4_7_0;
  assign ctb[7] = pp_4_7_1;
  assign cta[8] = pp_4_8_0;
  assign ctb[8] = pp_4_8_1;
  assign cta[9] = pp_4_9_0;
  assign ctb[9] = pp_4_9_1;
  assign cta[10] = pp_4_10_0;
  assign ctb[10] = pp_4_10_1;
  assign cta[11] = pp_4_11_0;
  assign ctb[11] = pp_4_11_1;
  assign cta[12] = pp_4_12_0;
  assign ctb[12] = pp_4_12_1;
  assign cta[13] = pp_4_13_0;
  assign ctb[13] = pp_4_13_1;
  assign cta[14] = pp_4_14_0;
  assign ctb[14] = pp_4_14_1;
  assign cta[15] = pp_4_15_0;
  assign ctb[15] = pp_4_15_1;
  assign cta[16] = pp_4_16_0;
  assign ctb[16] = pp_4_16_1;
  assign cta[17] = pp_4_17_0;
  assign ctb[17] = pp_4_17_1;
  assign cta[18] = pp_4_18_0;
  assign ctb[18] = pp_4_18_1;
  assign cta[19] = pp_4_19_0;
  assign ctb[19] = pp_4_19_1;
  assign cta[20] = pp_4_20_0;
  assign ctb[20] = pp_4_20_1;
  assign cta[21] = pp_4_21_0;
  assign ctb[21] = pp_4_21_1;
  assign cta[22] = pp_4_22_0;
  assign ctb[22] = pp_4_22_1;
  assign cta[23] = pp_4_23_0;
  assign ctb[23] = pp_4_23_1;
  assign cta[24] = pp_4_24_0;
  assign ctb[24] = pp_4_24_1;
  assign cta[25] = pp_4_25_0;
  assign ctb[25] = pp_4_25_1;
  assign cta[26] = pp_4_26_0;
  assign ctb[26] = pp_4_26_1;
  assign cta[27] = pp_4_27_0;
  assign ctb[27] = pp_4_27_1;
  assign cta[28] = pp_4_28_0;
  assign ctb[28] = pp_4_28_1;
  assign cta[29] = pp_4_29_0;
  assign ctb[29] = pp_4_29_1;
  assign cta[30] = pp_4_30_0;
  assign ctb[30] = pp_4_30_1;
  assign cta[31] = pp_4_31_0;
  assign ctb[31] = pp_4_31_1;
  assign product[31:0] = cts;
endmodule
