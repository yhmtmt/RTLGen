module MG_CPA(
  input [62:0] a,
  input [62:0] b,
  output [62:0] sum,
  output cout
);

  wire p_0_0;
  wire g_0_0;
 assign p_0_0 = a[0] ^ b[0];
 assign g_0_0 = a[0] & b[0];
  wire p_1_1;
  wire g_1_1;
 assign p_1_1 = a[1] ^ b[1];
 assign g_1_1 = a[1] & b[1];
  wire p_1_0;
  wire g_1_0;
  wire p_2_2;
  wire g_2_2;
 assign p_2_2 = a[2] ^ b[2];
 assign g_2_2 = a[2] & b[2];
  wire p_2_0;
  wire g_2_0;
  wire p_2_1;
  wire g_2_1;
  wire p_3_3;
  wire g_3_3;
 assign p_3_3 = a[3] ^ b[3];
 assign g_3_3 = a[3] & b[3];
  wire p_3_0;
  wire g_3_0;
  wire p_3_1;
  wire g_3_1;
  wire p_3_2;
  wire g_3_2;
  wire p_4_4;
  wire g_4_4;
 assign p_4_4 = a[4] ^ b[4];
 assign g_4_4 = a[4] & b[4];
  wire p_4_0;
  wire g_4_0;
  wire p_4_1;
  wire g_4_1;
  wire p_4_2;
  wire g_4_2;
  wire p_4_3;
  wire g_4_3;
  wire p_5_5;
  wire g_5_5;
 assign p_5_5 = a[5] ^ b[5];
 assign g_5_5 = a[5] & b[5];
  wire p_5_0;
  wire g_5_0;
  wire p_5_1;
  wire g_5_1;
  wire p_5_2;
  wire g_5_2;
  wire p_5_3;
  wire g_5_3;
  wire p_5_4;
  wire g_5_4;
  wire p_6_6;
  wire g_6_6;
 assign p_6_6 = a[6] ^ b[6];
 assign g_6_6 = a[6] & b[6];
  wire p_6_0;
  wire g_6_0;
  wire p_6_1;
  wire g_6_1;
  wire p_6_2;
  wire g_6_2;
  wire p_6_3;
  wire g_6_3;
  wire p_6_4;
  wire g_6_4;
  wire p_6_5;
  wire g_6_5;
  wire p_7_7;
  wire g_7_7;
 assign p_7_7 = a[7] ^ b[7];
 assign g_7_7 = a[7] & b[7];
  wire p_7_0;
  wire g_7_0;
  wire p_7_1;
  wire g_7_1;
  wire p_7_2;
  wire g_7_2;
  wire p_7_3;
  wire g_7_3;
  wire p_7_4;
  wire g_7_4;
  wire p_7_5;
  wire g_7_5;
  wire p_7_6;
  wire g_7_6;
  wire p_8_8;
  wire g_8_8;
 assign p_8_8 = a[8] ^ b[8];
 assign g_8_8 = a[8] & b[8];
  wire p_8_0;
  wire g_8_0;
  wire p_8_1;
  wire g_8_1;
  wire p_8_2;
  wire g_8_2;
  wire p_8_3;
  wire g_8_3;
  wire p_8_4;
  wire g_8_4;
  wire p_8_5;
  wire g_8_5;
  wire p_8_6;
  wire g_8_6;
  wire p_8_7;
  wire g_8_7;
  wire p_9_9;
  wire g_9_9;
 assign p_9_9 = a[9] ^ b[9];
 assign g_9_9 = a[9] & b[9];
  wire p_9_0;
  wire g_9_0;
  wire p_9_1;
  wire g_9_1;
  wire p_9_2;
  wire g_9_2;
  wire p_9_3;
  wire g_9_3;
  wire p_9_4;
  wire g_9_4;
  wire p_9_5;
  wire g_9_5;
  wire p_9_6;
  wire g_9_6;
  wire p_9_7;
  wire g_9_7;
  wire p_9_8;
  wire g_9_8;
  wire p_10_10;
  wire g_10_10;
 assign p_10_10 = a[10] ^ b[10];
 assign g_10_10 = a[10] & b[10];
  wire p_10_0;
  wire g_10_0;
  wire p_10_1;
  wire g_10_1;
  wire p_10_2;
  wire g_10_2;
  wire p_10_3;
  wire g_10_3;
  wire p_10_4;
  wire g_10_4;
  wire p_10_5;
  wire g_10_5;
  wire p_10_6;
  wire g_10_6;
  wire p_10_7;
  wire g_10_7;
  wire p_10_8;
  wire g_10_8;
  wire p_10_9;
  wire g_10_9;
  wire p_11_11;
  wire g_11_11;
 assign p_11_11 = a[11] ^ b[11];
 assign g_11_11 = a[11] & b[11];
  wire p_11_0;
  wire g_11_0;
  wire p_11_1;
  wire g_11_1;
  wire p_11_2;
  wire g_11_2;
  wire p_11_3;
  wire g_11_3;
  wire p_11_4;
  wire g_11_4;
  wire p_11_5;
  wire g_11_5;
  wire p_11_6;
  wire g_11_6;
  wire p_11_7;
  wire g_11_7;
  wire p_11_8;
  wire g_11_8;
  wire p_11_9;
  wire g_11_9;
  wire p_11_10;
  wire g_11_10;
  wire p_12_12;
  wire g_12_12;
 assign p_12_12 = a[12] ^ b[12];
 assign g_12_12 = a[12] & b[12];
  wire p_12_0;
  wire g_12_0;
  wire p_12_1;
  wire g_12_1;
  wire p_12_2;
  wire g_12_2;
  wire p_12_3;
  wire g_12_3;
  wire p_12_4;
  wire g_12_4;
  wire p_12_5;
  wire g_12_5;
  wire p_12_6;
  wire g_12_6;
  wire p_12_7;
  wire g_12_7;
  wire p_12_8;
  wire g_12_8;
  wire p_12_9;
  wire g_12_9;
  wire p_12_10;
  wire g_12_10;
  wire p_12_11;
  wire g_12_11;
  wire p_13_13;
  wire g_13_13;
 assign p_13_13 = a[13] ^ b[13];
 assign g_13_13 = a[13] & b[13];
  wire p_13_0;
  wire g_13_0;
  wire p_13_1;
  wire g_13_1;
  wire p_13_2;
  wire g_13_2;
  wire p_13_3;
  wire g_13_3;
  wire p_13_4;
  wire g_13_4;
  wire p_13_5;
  wire g_13_5;
  wire p_13_6;
  wire g_13_6;
  wire p_13_7;
  wire g_13_7;
  wire p_13_8;
  wire g_13_8;
  wire p_13_9;
  wire g_13_9;
  wire p_13_10;
  wire g_13_10;
  wire p_13_11;
  wire g_13_11;
  wire p_13_12;
  wire g_13_12;
  wire p_14_14;
  wire g_14_14;
 assign p_14_14 = a[14] ^ b[14];
 assign g_14_14 = a[14] & b[14];
  wire p_14_0;
  wire g_14_0;
  wire p_14_1;
  wire g_14_1;
  wire p_14_2;
  wire g_14_2;
  wire p_14_3;
  wire g_14_3;
  wire p_14_4;
  wire g_14_4;
  wire p_14_5;
  wire g_14_5;
  wire p_14_6;
  wire g_14_6;
  wire p_14_7;
  wire g_14_7;
  wire p_14_8;
  wire g_14_8;
  wire p_14_9;
  wire g_14_9;
  wire p_14_10;
  wire g_14_10;
  wire p_14_11;
  wire g_14_11;
  wire p_14_12;
  wire g_14_12;
  wire p_14_13;
  wire g_14_13;
  wire p_15_15;
  wire g_15_15;
 assign p_15_15 = a[15] ^ b[15];
 assign g_15_15 = a[15] & b[15];
  wire p_15_0;
  wire g_15_0;
  wire p_15_1;
  wire g_15_1;
  wire p_15_2;
  wire g_15_2;
  wire p_15_3;
  wire g_15_3;
  wire p_15_4;
  wire g_15_4;
  wire p_15_5;
  wire g_15_5;
  wire p_15_6;
  wire g_15_6;
  wire p_15_7;
  wire g_15_7;
  wire p_15_8;
  wire g_15_8;
  wire p_15_9;
  wire g_15_9;
  wire p_15_10;
  wire g_15_10;
  wire p_15_11;
  wire g_15_11;
  wire p_15_12;
  wire g_15_12;
  wire p_15_13;
  wire g_15_13;
  wire p_15_14;
  wire g_15_14;
  wire p_16_16;
  wire g_16_16;
 assign p_16_16 = a[16] ^ b[16];
 assign g_16_16 = a[16] & b[16];
  wire p_16_0;
  wire g_16_0;
  wire p_16_1;
  wire g_16_1;
  wire p_16_2;
  wire g_16_2;
  wire p_16_3;
  wire g_16_3;
  wire p_16_4;
  wire g_16_4;
  wire p_16_5;
  wire g_16_5;
  wire p_16_6;
  wire g_16_6;
  wire p_16_7;
  wire g_16_7;
  wire p_16_8;
  wire g_16_8;
  wire p_16_9;
  wire g_16_9;
  wire p_16_10;
  wire g_16_10;
  wire p_16_11;
  wire g_16_11;
  wire p_16_12;
  wire g_16_12;
  wire p_16_13;
  wire g_16_13;
  wire p_16_14;
  wire g_16_14;
  wire p_16_15;
  wire g_16_15;
  wire p_17_17;
  wire g_17_17;
 assign p_17_17 = a[17] ^ b[17];
 assign g_17_17 = a[17] & b[17];
  wire p_17_0;
  wire g_17_0;
  wire p_17_1;
  wire g_17_1;
  wire p_17_2;
  wire g_17_2;
  wire p_17_3;
  wire g_17_3;
  wire p_17_4;
  wire g_17_4;
  wire p_17_5;
  wire g_17_5;
  wire p_17_6;
  wire g_17_6;
  wire p_17_7;
  wire g_17_7;
  wire p_17_8;
  wire g_17_8;
  wire p_17_9;
  wire g_17_9;
  wire p_17_10;
  wire g_17_10;
  wire p_17_11;
  wire g_17_11;
  wire p_17_12;
  wire g_17_12;
  wire p_17_13;
  wire g_17_13;
  wire p_17_14;
  wire g_17_14;
  wire p_17_15;
  wire g_17_15;
  wire p_17_16;
  wire g_17_16;
  wire p_18_18;
  wire g_18_18;
 assign p_18_18 = a[18] ^ b[18];
 assign g_18_18 = a[18] & b[18];
  wire p_18_0;
  wire g_18_0;
  wire p_18_1;
  wire g_18_1;
  wire p_18_2;
  wire g_18_2;
  wire p_18_3;
  wire g_18_3;
  wire p_18_4;
  wire g_18_4;
  wire p_18_5;
  wire g_18_5;
  wire p_18_6;
  wire g_18_6;
  wire p_18_7;
  wire g_18_7;
  wire p_18_8;
  wire g_18_8;
  wire p_18_9;
  wire g_18_9;
  wire p_18_10;
  wire g_18_10;
  wire p_18_11;
  wire g_18_11;
  wire p_18_12;
  wire g_18_12;
  wire p_18_13;
  wire g_18_13;
  wire p_18_14;
  wire g_18_14;
  wire p_18_15;
  wire g_18_15;
  wire p_18_16;
  wire g_18_16;
  wire p_18_17;
  wire g_18_17;
  wire p_19_19;
  wire g_19_19;
 assign p_19_19 = a[19] ^ b[19];
 assign g_19_19 = a[19] & b[19];
  wire p_19_0;
  wire g_19_0;
  wire p_19_1;
  wire g_19_1;
  wire p_19_2;
  wire g_19_2;
  wire p_19_3;
  wire g_19_3;
  wire p_19_4;
  wire g_19_4;
  wire p_19_5;
  wire g_19_5;
  wire p_19_6;
  wire g_19_6;
  wire p_19_7;
  wire g_19_7;
  wire p_19_8;
  wire g_19_8;
  wire p_19_9;
  wire g_19_9;
  wire p_19_10;
  wire g_19_10;
  wire p_19_11;
  wire g_19_11;
  wire p_19_12;
  wire g_19_12;
  wire p_19_13;
  wire g_19_13;
  wire p_19_14;
  wire g_19_14;
  wire p_19_15;
  wire g_19_15;
  wire p_19_16;
  wire g_19_16;
  wire p_19_17;
  wire g_19_17;
  wire p_19_18;
  wire g_19_18;
  wire p_20_20;
  wire g_20_20;
 assign p_20_20 = a[20] ^ b[20];
 assign g_20_20 = a[20] & b[20];
  wire p_20_0;
  wire g_20_0;
  wire p_20_1;
  wire g_20_1;
  wire p_20_2;
  wire g_20_2;
  wire p_20_3;
  wire g_20_3;
  wire p_20_4;
  wire g_20_4;
  wire p_20_5;
  wire g_20_5;
  wire p_20_6;
  wire g_20_6;
  wire p_20_7;
  wire g_20_7;
  wire p_20_8;
  wire g_20_8;
  wire p_20_9;
  wire g_20_9;
  wire p_20_10;
  wire g_20_10;
  wire p_20_11;
  wire g_20_11;
  wire p_20_12;
  wire g_20_12;
  wire p_20_13;
  wire g_20_13;
  wire p_20_14;
  wire g_20_14;
  wire p_20_15;
  wire g_20_15;
  wire p_20_16;
  wire g_20_16;
  wire p_20_17;
  wire g_20_17;
  wire p_20_18;
  wire g_20_18;
  wire p_20_19;
  wire g_20_19;
  wire p_21_21;
  wire g_21_21;
 assign p_21_21 = a[21] ^ b[21];
 assign g_21_21 = a[21] & b[21];
  wire p_21_0;
  wire g_21_0;
  wire p_21_1;
  wire g_21_1;
  wire p_21_2;
  wire g_21_2;
  wire p_21_3;
  wire g_21_3;
  wire p_21_4;
  wire g_21_4;
  wire p_21_5;
  wire g_21_5;
  wire p_21_6;
  wire g_21_6;
  wire p_21_7;
  wire g_21_7;
  wire p_21_8;
  wire g_21_8;
  wire p_21_9;
  wire g_21_9;
  wire p_21_10;
  wire g_21_10;
  wire p_21_11;
  wire g_21_11;
  wire p_21_12;
  wire g_21_12;
  wire p_21_13;
  wire g_21_13;
  wire p_21_14;
  wire g_21_14;
  wire p_21_15;
  wire g_21_15;
  wire p_21_16;
  wire g_21_16;
  wire p_21_17;
  wire g_21_17;
  wire p_21_18;
  wire g_21_18;
  wire p_21_19;
  wire g_21_19;
  wire p_21_20;
  wire g_21_20;
  wire p_22_22;
  wire g_22_22;
 assign p_22_22 = a[22] ^ b[22];
 assign g_22_22 = a[22] & b[22];
  wire p_22_0;
  wire g_22_0;
  wire p_22_1;
  wire g_22_1;
  wire p_22_2;
  wire g_22_2;
  wire p_22_3;
  wire g_22_3;
  wire p_22_4;
  wire g_22_4;
  wire p_22_5;
  wire g_22_5;
  wire p_22_6;
  wire g_22_6;
  wire p_22_7;
  wire g_22_7;
  wire p_22_8;
  wire g_22_8;
  wire p_22_9;
  wire g_22_9;
  wire p_22_10;
  wire g_22_10;
  wire p_22_11;
  wire g_22_11;
  wire p_22_12;
  wire g_22_12;
  wire p_22_13;
  wire g_22_13;
  wire p_22_14;
  wire g_22_14;
  wire p_22_15;
  wire g_22_15;
  wire p_22_16;
  wire g_22_16;
  wire p_22_17;
  wire g_22_17;
  wire p_22_18;
  wire g_22_18;
  wire p_22_19;
  wire g_22_19;
  wire p_22_20;
  wire g_22_20;
  wire p_22_21;
  wire g_22_21;
  wire p_23_23;
  wire g_23_23;
 assign p_23_23 = a[23] ^ b[23];
 assign g_23_23 = a[23] & b[23];
  wire p_23_0;
  wire g_23_0;
  wire p_23_1;
  wire g_23_1;
  wire p_23_2;
  wire g_23_2;
  wire p_23_3;
  wire g_23_3;
  wire p_23_4;
  wire g_23_4;
  wire p_23_5;
  wire g_23_5;
  wire p_23_6;
  wire g_23_6;
  wire p_23_7;
  wire g_23_7;
  wire p_23_8;
  wire g_23_8;
  wire p_23_9;
  wire g_23_9;
  wire p_23_10;
  wire g_23_10;
  wire p_23_11;
  wire g_23_11;
  wire p_23_12;
  wire g_23_12;
  wire p_23_13;
  wire g_23_13;
  wire p_23_14;
  wire g_23_14;
  wire p_23_15;
  wire g_23_15;
  wire p_23_16;
  wire g_23_16;
  wire p_23_17;
  wire g_23_17;
  wire p_23_18;
  wire g_23_18;
  wire p_23_19;
  wire g_23_19;
  wire p_23_20;
  wire g_23_20;
  wire p_23_21;
  wire g_23_21;
  wire p_23_22;
  wire g_23_22;
  wire p_24_24;
  wire g_24_24;
 assign p_24_24 = a[24] ^ b[24];
 assign g_24_24 = a[24] & b[24];
  wire p_24_0;
  wire g_24_0;
  wire p_24_1;
  wire g_24_1;
  wire p_24_2;
  wire g_24_2;
  wire p_24_3;
  wire g_24_3;
  wire p_24_4;
  wire g_24_4;
  wire p_24_5;
  wire g_24_5;
  wire p_24_6;
  wire g_24_6;
  wire p_24_7;
  wire g_24_7;
  wire p_24_8;
  wire g_24_8;
  wire p_24_9;
  wire g_24_9;
  wire p_24_10;
  wire g_24_10;
  wire p_24_11;
  wire g_24_11;
  wire p_24_12;
  wire g_24_12;
  wire p_24_13;
  wire g_24_13;
  wire p_24_14;
  wire g_24_14;
  wire p_24_15;
  wire g_24_15;
  wire p_24_16;
  wire g_24_16;
  wire p_24_17;
  wire g_24_17;
  wire p_24_18;
  wire g_24_18;
  wire p_24_19;
  wire g_24_19;
  wire p_24_20;
  wire g_24_20;
  wire p_24_21;
  wire g_24_21;
  wire p_24_22;
  wire g_24_22;
  wire p_24_23;
  wire g_24_23;
  wire p_25_25;
  wire g_25_25;
 assign p_25_25 = a[25] ^ b[25];
 assign g_25_25 = a[25] & b[25];
  wire p_25_0;
  wire g_25_0;
  wire p_25_1;
  wire g_25_1;
  wire p_25_2;
  wire g_25_2;
  wire p_25_3;
  wire g_25_3;
  wire p_25_4;
  wire g_25_4;
  wire p_25_5;
  wire g_25_5;
  wire p_25_6;
  wire g_25_6;
  wire p_25_7;
  wire g_25_7;
  wire p_25_8;
  wire g_25_8;
  wire p_25_9;
  wire g_25_9;
  wire p_25_10;
  wire g_25_10;
  wire p_25_11;
  wire g_25_11;
  wire p_25_12;
  wire g_25_12;
  wire p_25_13;
  wire g_25_13;
  wire p_25_14;
  wire g_25_14;
  wire p_25_15;
  wire g_25_15;
  wire p_25_16;
  wire g_25_16;
  wire p_25_17;
  wire g_25_17;
  wire p_25_18;
  wire g_25_18;
  wire p_25_19;
  wire g_25_19;
  wire p_25_20;
  wire g_25_20;
  wire p_25_21;
  wire g_25_21;
  wire p_25_22;
  wire g_25_22;
  wire p_25_23;
  wire g_25_23;
  wire p_25_24;
  wire g_25_24;
  wire p_26_26;
  wire g_26_26;
 assign p_26_26 = a[26] ^ b[26];
 assign g_26_26 = a[26] & b[26];
  wire p_26_0;
  wire g_26_0;
  wire p_26_1;
  wire g_26_1;
  wire p_26_2;
  wire g_26_2;
  wire p_26_3;
  wire g_26_3;
  wire p_26_4;
  wire g_26_4;
  wire p_26_5;
  wire g_26_5;
  wire p_26_6;
  wire g_26_6;
  wire p_26_7;
  wire g_26_7;
  wire p_26_8;
  wire g_26_8;
  wire p_26_9;
  wire g_26_9;
  wire p_26_10;
  wire g_26_10;
  wire p_26_11;
  wire g_26_11;
  wire p_26_12;
  wire g_26_12;
  wire p_26_13;
  wire g_26_13;
  wire p_26_14;
  wire g_26_14;
  wire p_26_15;
  wire g_26_15;
  wire p_26_16;
  wire g_26_16;
  wire p_26_17;
  wire g_26_17;
  wire p_26_18;
  wire g_26_18;
  wire p_26_19;
  wire g_26_19;
  wire p_26_20;
  wire g_26_20;
  wire p_26_21;
  wire g_26_21;
  wire p_26_22;
  wire g_26_22;
  wire p_26_23;
  wire g_26_23;
  wire p_26_24;
  wire g_26_24;
  wire p_26_25;
  wire g_26_25;
  wire p_27_27;
  wire g_27_27;
 assign p_27_27 = a[27] ^ b[27];
 assign g_27_27 = a[27] & b[27];
  wire p_27_0;
  wire g_27_0;
  wire p_27_1;
  wire g_27_1;
  wire p_27_2;
  wire g_27_2;
  wire p_27_3;
  wire g_27_3;
  wire p_27_4;
  wire g_27_4;
  wire p_27_5;
  wire g_27_5;
  wire p_27_6;
  wire g_27_6;
  wire p_27_7;
  wire g_27_7;
  wire p_27_8;
  wire g_27_8;
  wire p_27_9;
  wire g_27_9;
  wire p_27_10;
  wire g_27_10;
  wire p_27_11;
  wire g_27_11;
  wire p_27_12;
  wire g_27_12;
  wire p_27_13;
  wire g_27_13;
  wire p_27_14;
  wire g_27_14;
  wire p_27_15;
  wire g_27_15;
  wire p_27_16;
  wire g_27_16;
  wire p_27_17;
  wire g_27_17;
  wire p_27_18;
  wire g_27_18;
  wire p_27_19;
  wire g_27_19;
  wire p_27_20;
  wire g_27_20;
  wire p_27_21;
  wire g_27_21;
  wire p_27_22;
  wire g_27_22;
  wire p_27_23;
  wire g_27_23;
  wire p_27_24;
  wire g_27_24;
  wire p_27_25;
  wire g_27_25;
  wire p_27_26;
  wire g_27_26;
  wire p_28_28;
  wire g_28_28;
 assign p_28_28 = a[28] ^ b[28];
 assign g_28_28 = a[28] & b[28];
  wire p_28_0;
  wire g_28_0;
  wire p_28_1;
  wire g_28_1;
  wire p_28_2;
  wire g_28_2;
  wire p_28_3;
  wire g_28_3;
  wire p_28_4;
  wire g_28_4;
  wire p_28_5;
  wire g_28_5;
  wire p_28_6;
  wire g_28_6;
  wire p_28_7;
  wire g_28_7;
  wire p_28_8;
  wire g_28_8;
  wire p_28_9;
  wire g_28_9;
  wire p_28_10;
  wire g_28_10;
  wire p_28_11;
  wire g_28_11;
  wire p_28_12;
  wire g_28_12;
  wire p_28_13;
  wire g_28_13;
  wire p_28_14;
  wire g_28_14;
  wire p_28_15;
  wire g_28_15;
  wire p_28_16;
  wire g_28_16;
  wire p_28_17;
  wire g_28_17;
  wire p_28_18;
  wire g_28_18;
  wire p_28_19;
  wire g_28_19;
  wire p_28_20;
  wire g_28_20;
  wire p_28_21;
  wire g_28_21;
  wire p_28_22;
  wire g_28_22;
  wire p_28_23;
  wire g_28_23;
  wire p_28_24;
  wire g_28_24;
  wire p_28_25;
  wire g_28_25;
  wire p_28_26;
  wire g_28_26;
  wire p_28_27;
  wire g_28_27;
  wire p_29_29;
  wire g_29_29;
 assign p_29_29 = a[29] ^ b[29];
 assign g_29_29 = a[29] & b[29];
  wire p_29_0;
  wire g_29_0;
  wire p_29_1;
  wire g_29_1;
  wire p_29_2;
  wire g_29_2;
  wire p_29_3;
  wire g_29_3;
  wire p_29_4;
  wire g_29_4;
  wire p_29_5;
  wire g_29_5;
  wire p_29_6;
  wire g_29_6;
  wire p_29_7;
  wire g_29_7;
  wire p_29_8;
  wire g_29_8;
  wire p_29_9;
  wire g_29_9;
  wire p_29_10;
  wire g_29_10;
  wire p_29_11;
  wire g_29_11;
  wire p_29_12;
  wire g_29_12;
  wire p_29_13;
  wire g_29_13;
  wire p_29_14;
  wire g_29_14;
  wire p_29_15;
  wire g_29_15;
  wire p_29_16;
  wire g_29_16;
  wire p_29_17;
  wire g_29_17;
  wire p_29_18;
  wire g_29_18;
  wire p_29_19;
  wire g_29_19;
  wire p_29_20;
  wire g_29_20;
  wire p_29_21;
  wire g_29_21;
  wire p_29_22;
  wire g_29_22;
  wire p_29_23;
  wire g_29_23;
  wire p_29_24;
  wire g_29_24;
  wire p_29_25;
  wire g_29_25;
  wire p_29_26;
  wire g_29_26;
  wire p_29_27;
  wire g_29_27;
  wire p_29_28;
  wire g_29_28;
  wire p_30_30;
  wire g_30_30;
 assign p_30_30 = a[30] ^ b[30];
 assign g_30_30 = a[30] & b[30];
  wire p_30_0;
  wire g_30_0;
  wire p_30_1;
  wire g_30_1;
  wire p_30_2;
  wire g_30_2;
  wire p_30_3;
  wire g_30_3;
  wire p_30_4;
  wire g_30_4;
  wire p_30_5;
  wire g_30_5;
  wire p_30_6;
  wire g_30_6;
  wire p_30_7;
  wire g_30_7;
  wire p_30_8;
  wire g_30_8;
  wire p_30_9;
  wire g_30_9;
  wire p_30_10;
  wire g_30_10;
  wire p_30_11;
  wire g_30_11;
  wire p_30_12;
  wire g_30_12;
  wire p_30_13;
  wire g_30_13;
  wire p_30_14;
  wire g_30_14;
  wire p_30_15;
  wire g_30_15;
  wire p_30_16;
  wire g_30_16;
  wire p_30_17;
  wire g_30_17;
  wire p_30_18;
  wire g_30_18;
  wire p_30_19;
  wire g_30_19;
  wire p_30_20;
  wire g_30_20;
  wire p_30_21;
  wire g_30_21;
  wire p_30_22;
  wire g_30_22;
  wire p_30_23;
  wire g_30_23;
  wire p_30_24;
  wire g_30_24;
  wire p_30_25;
  wire g_30_25;
  wire p_30_26;
  wire g_30_26;
  wire p_30_27;
  wire g_30_27;
  wire p_30_28;
  wire g_30_28;
  wire p_30_29;
  wire g_30_29;
  wire p_31_31;
  wire g_31_31;
 assign p_31_31 = a[31] ^ b[31];
 assign g_31_31 = a[31] & b[31];
  wire p_31_0;
  wire g_31_0;
  wire p_31_1;
  wire g_31_1;
  wire p_31_2;
  wire g_31_2;
  wire p_31_3;
  wire g_31_3;
  wire p_31_4;
  wire g_31_4;
  wire p_31_5;
  wire g_31_5;
  wire p_31_6;
  wire g_31_6;
  wire p_31_7;
  wire g_31_7;
  wire p_31_8;
  wire g_31_8;
  wire p_31_9;
  wire g_31_9;
  wire p_31_10;
  wire g_31_10;
  wire p_31_11;
  wire g_31_11;
  wire p_31_12;
  wire g_31_12;
  wire p_31_13;
  wire g_31_13;
  wire p_31_14;
  wire g_31_14;
  wire p_31_15;
  wire g_31_15;
  wire p_31_16;
  wire g_31_16;
  wire p_31_17;
  wire g_31_17;
  wire p_31_18;
  wire g_31_18;
  wire p_31_19;
  wire g_31_19;
  wire p_31_20;
  wire g_31_20;
  wire p_31_21;
  wire g_31_21;
  wire p_31_22;
  wire g_31_22;
  wire p_31_23;
  wire g_31_23;
  wire p_31_24;
  wire g_31_24;
  wire p_31_25;
  wire g_31_25;
  wire p_31_26;
  wire g_31_26;
  wire p_31_27;
  wire g_31_27;
  wire p_31_28;
  wire g_31_28;
  wire p_31_29;
  wire g_31_29;
  wire p_31_30;
  wire g_31_30;
  wire p_32_32;
  wire g_32_32;
 assign p_32_32 = a[32] ^ b[32];
 assign g_32_32 = a[32] & b[32];
  wire p_32_0;
  wire g_32_0;
  wire p_32_1;
  wire g_32_1;
  wire p_32_2;
  wire g_32_2;
  wire p_32_3;
  wire g_32_3;
  wire p_32_4;
  wire g_32_4;
  wire p_32_5;
  wire g_32_5;
  wire p_32_6;
  wire g_32_6;
  wire p_32_7;
  wire g_32_7;
  wire p_32_8;
  wire g_32_8;
  wire p_32_9;
  wire g_32_9;
  wire p_32_10;
  wire g_32_10;
  wire p_32_11;
  wire g_32_11;
  wire p_32_12;
  wire g_32_12;
  wire p_32_13;
  wire g_32_13;
  wire p_32_14;
  wire g_32_14;
  wire p_32_15;
  wire g_32_15;
  wire p_32_16;
  wire g_32_16;
  wire p_32_17;
  wire g_32_17;
  wire p_32_18;
  wire g_32_18;
  wire p_32_19;
  wire g_32_19;
  wire p_32_20;
  wire g_32_20;
  wire p_32_21;
  wire g_32_21;
  wire p_32_22;
  wire g_32_22;
  wire p_32_23;
  wire g_32_23;
  wire p_32_24;
  wire g_32_24;
  wire p_32_25;
  wire g_32_25;
  wire p_32_26;
  wire g_32_26;
  wire p_32_27;
  wire g_32_27;
  wire p_32_28;
  wire g_32_28;
  wire p_32_29;
  wire g_32_29;
  wire p_32_30;
  wire g_32_30;
  wire p_32_31;
  wire g_32_31;
  wire p_33_33;
  wire g_33_33;
 assign p_33_33 = a[33] ^ b[33];
 assign g_33_33 = a[33] & b[33];
  wire p_33_0;
  wire g_33_0;
  wire p_33_1;
  wire g_33_1;
  wire p_33_2;
  wire g_33_2;
  wire p_33_3;
  wire g_33_3;
  wire p_33_4;
  wire g_33_4;
  wire p_33_5;
  wire g_33_5;
  wire p_33_6;
  wire g_33_6;
  wire p_33_7;
  wire g_33_7;
  wire p_33_8;
  wire g_33_8;
  wire p_33_9;
  wire g_33_9;
  wire p_33_10;
  wire g_33_10;
  wire p_33_11;
  wire g_33_11;
  wire p_33_12;
  wire g_33_12;
  wire p_33_13;
  wire g_33_13;
  wire p_33_14;
  wire g_33_14;
  wire p_33_15;
  wire g_33_15;
  wire p_33_16;
  wire g_33_16;
  wire p_33_17;
  wire g_33_17;
  wire p_33_18;
  wire g_33_18;
  wire p_33_19;
  wire g_33_19;
  wire p_33_20;
  wire g_33_20;
  wire p_33_21;
  wire g_33_21;
  wire p_33_22;
  wire g_33_22;
  wire p_33_23;
  wire g_33_23;
  wire p_33_24;
  wire g_33_24;
  wire p_33_25;
  wire g_33_25;
  wire p_33_26;
  wire g_33_26;
  wire p_33_27;
  wire g_33_27;
  wire p_33_28;
  wire g_33_28;
  wire p_33_29;
  wire g_33_29;
  wire p_33_30;
  wire g_33_30;
  wire p_33_31;
  wire g_33_31;
  wire p_33_32;
  wire g_33_32;
  wire p_34_34;
  wire g_34_34;
 assign p_34_34 = a[34] ^ b[34];
 assign g_34_34 = a[34] & b[34];
  wire p_34_0;
  wire g_34_0;
  wire p_34_1;
  wire g_34_1;
  wire p_34_2;
  wire g_34_2;
  wire p_34_3;
  wire g_34_3;
  wire p_34_4;
  wire g_34_4;
  wire p_34_5;
  wire g_34_5;
  wire p_34_6;
  wire g_34_6;
  wire p_34_7;
  wire g_34_7;
  wire p_34_8;
  wire g_34_8;
  wire p_34_9;
  wire g_34_9;
  wire p_34_10;
  wire g_34_10;
  wire p_34_11;
  wire g_34_11;
  wire p_34_12;
  wire g_34_12;
  wire p_34_13;
  wire g_34_13;
  wire p_34_14;
  wire g_34_14;
  wire p_34_15;
  wire g_34_15;
  wire p_34_16;
  wire g_34_16;
  wire p_34_17;
  wire g_34_17;
  wire p_34_18;
  wire g_34_18;
  wire p_34_19;
  wire g_34_19;
  wire p_34_20;
  wire g_34_20;
  wire p_34_21;
  wire g_34_21;
  wire p_34_22;
  wire g_34_22;
  wire p_34_23;
  wire g_34_23;
  wire p_34_24;
  wire g_34_24;
  wire p_34_25;
  wire g_34_25;
  wire p_34_26;
  wire g_34_26;
  wire p_34_27;
  wire g_34_27;
  wire p_34_28;
  wire g_34_28;
  wire p_34_29;
  wire g_34_29;
  wire p_34_30;
  wire g_34_30;
  wire p_34_31;
  wire g_34_31;
  wire p_34_32;
  wire g_34_32;
  wire p_34_33;
  wire g_34_33;
  wire p_35_35;
  wire g_35_35;
 assign p_35_35 = a[35] ^ b[35];
 assign g_35_35 = a[35] & b[35];
  wire p_35_0;
  wire g_35_0;
  wire p_35_1;
  wire g_35_1;
  wire p_35_2;
  wire g_35_2;
  wire p_35_3;
  wire g_35_3;
  wire p_35_4;
  wire g_35_4;
  wire p_35_5;
  wire g_35_5;
  wire p_35_6;
  wire g_35_6;
  wire p_35_7;
  wire g_35_7;
  wire p_35_8;
  wire g_35_8;
  wire p_35_9;
  wire g_35_9;
  wire p_35_10;
  wire g_35_10;
  wire p_35_11;
  wire g_35_11;
  wire p_35_12;
  wire g_35_12;
  wire p_35_13;
  wire g_35_13;
  wire p_35_14;
  wire g_35_14;
  wire p_35_15;
  wire g_35_15;
  wire p_35_16;
  wire g_35_16;
  wire p_35_17;
  wire g_35_17;
  wire p_35_18;
  wire g_35_18;
  wire p_35_19;
  wire g_35_19;
  wire p_35_20;
  wire g_35_20;
  wire p_35_21;
  wire g_35_21;
  wire p_35_22;
  wire g_35_22;
  wire p_35_23;
  wire g_35_23;
  wire p_35_24;
  wire g_35_24;
  wire p_35_25;
  wire g_35_25;
  wire p_35_26;
  wire g_35_26;
  wire p_35_27;
  wire g_35_27;
  wire p_35_28;
  wire g_35_28;
  wire p_35_29;
  wire g_35_29;
  wire p_35_30;
  wire g_35_30;
  wire p_35_31;
  wire g_35_31;
  wire p_35_32;
  wire g_35_32;
  wire p_35_33;
  wire g_35_33;
  wire p_35_34;
  wire g_35_34;
  wire p_36_36;
  wire g_36_36;
 assign p_36_36 = a[36] ^ b[36];
 assign g_36_36 = a[36] & b[36];
  wire p_36_0;
  wire g_36_0;
  wire p_36_1;
  wire g_36_1;
  wire p_36_2;
  wire g_36_2;
  wire p_36_3;
  wire g_36_3;
  wire p_36_4;
  wire g_36_4;
  wire p_36_5;
  wire g_36_5;
  wire p_36_6;
  wire g_36_6;
  wire p_36_7;
  wire g_36_7;
  wire p_36_8;
  wire g_36_8;
  wire p_36_9;
  wire g_36_9;
  wire p_36_10;
  wire g_36_10;
  wire p_36_11;
  wire g_36_11;
  wire p_36_12;
  wire g_36_12;
  wire p_36_13;
  wire g_36_13;
  wire p_36_14;
  wire g_36_14;
  wire p_36_15;
  wire g_36_15;
  wire p_36_16;
  wire g_36_16;
  wire p_36_17;
  wire g_36_17;
  wire p_36_18;
  wire g_36_18;
  wire p_36_19;
  wire g_36_19;
  wire p_36_20;
  wire g_36_20;
  wire p_36_21;
  wire g_36_21;
  wire p_36_22;
  wire g_36_22;
  wire p_36_23;
  wire g_36_23;
  wire p_36_24;
  wire g_36_24;
  wire p_36_25;
  wire g_36_25;
  wire p_36_26;
  wire g_36_26;
  wire p_36_27;
  wire g_36_27;
  wire p_36_28;
  wire g_36_28;
  wire p_36_29;
  wire g_36_29;
  wire p_36_30;
  wire g_36_30;
  wire p_36_31;
  wire g_36_31;
  wire p_36_32;
  wire g_36_32;
  wire p_36_33;
  wire g_36_33;
  wire p_36_34;
  wire g_36_34;
  wire p_36_35;
  wire g_36_35;
  wire p_37_37;
  wire g_37_37;
 assign p_37_37 = a[37] ^ b[37];
 assign g_37_37 = a[37] & b[37];
  wire p_37_0;
  wire g_37_0;
  wire p_37_1;
  wire g_37_1;
  wire p_37_2;
  wire g_37_2;
  wire p_37_3;
  wire g_37_3;
  wire p_37_4;
  wire g_37_4;
  wire p_37_5;
  wire g_37_5;
  wire p_37_6;
  wire g_37_6;
  wire p_37_7;
  wire g_37_7;
  wire p_37_8;
  wire g_37_8;
  wire p_37_9;
  wire g_37_9;
  wire p_37_10;
  wire g_37_10;
  wire p_37_11;
  wire g_37_11;
  wire p_37_12;
  wire g_37_12;
  wire p_37_13;
  wire g_37_13;
  wire p_37_14;
  wire g_37_14;
  wire p_37_15;
  wire g_37_15;
  wire p_37_16;
  wire g_37_16;
  wire p_37_17;
  wire g_37_17;
  wire p_37_18;
  wire g_37_18;
  wire p_37_19;
  wire g_37_19;
  wire p_37_20;
  wire g_37_20;
  wire p_37_21;
  wire g_37_21;
  wire p_37_22;
  wire g_37_22;
  wire p_37_23;
  wire g_37_23;
  wire p_37_24;
  wire g_37_24;
  wire p_37_25;
  wire g_37_25;
  wire p_37_26;
  wire g_37_26;
  wire p_37_27;
  wire g_37_27;
  wire p_37_28;
  wire g_37_28;
  wire p_37_29;
  wire g_37_29;
  wire p_37_30;
  wire g_37_30;
  wire p_37_31;
  wire g_37_31;
  wire p_37_32;
  wire g_37_32;
  wire p_37_33;
  wire g_37_33;
  wire p_37_34;
  wire g_37_34;
  wire p_37_35;
  wire g_37_35;
  wire p_37_36;
  wire g_37_36;
  wire p_38_38;
  wire g_38_38;
 assign p_38_38 = a[38] ^ b[38];
 assign g_38_38 = a[38] & b[38];
  wire p_38_0;
  wire g_38_0;
  wire p_38_1;
  wire g_38_1;
  wire p_38_2;
  wire g_38_2;
  wire p_38_3;
  wire g_38_3;
  wire p_38_4;
  wire g_38_4;
  wire p_38_5;
  wire g_38_5;
  wire p_38_6;
  wire g_38_6;
  wire p_38_7;
  wire g_38_7;
  wire p_38_8;
  wire g_38_8;
  wire p_38_9;
  wire g_38_9;
  wire p_38_10;
  wire g_38_10;
  wire p_38_11;
  wire g_38_11;
  wire p_38_12;
  wire g_38_12;
  wire p_38_13;
  wire g_38_13;
  wire p_38_14;
  wire g_38_14;
  wire p_38_15;
  wire g_38_15;
  wire p_38_16;
  wire g_38_16;
  wire p_38_17;
  wire g_38_17;
  wire p_38_18;
  wire g_38_18;
  wire p_38_19;
  wire g_38_19;
  wire p_38_20;
  wire g_38_20;
  wire p_38_21;
  wire g_38_21;
  wire p_38_22;
  wire g_38_22;
  wire p_38_23;
  wire g_38_23;
  wire p_38_24;
  wire g_38_24;
  wire p_38_25;
  wire g_38_25;
  wire p_38_26;
  wire g_38_26;
  wire p_38_27;
  wire g_38_27;
  wire p_38_28;
  wire g_38_28;
  wire p_38_29;
  wire g_38_29;
  wire p_38_30;
  wire g_38_30;
  wire p_38_31;
  wire g_38_31;
  wire p_38_32;
  wire g_38_32;
  wire p_38_33;
  wire g_38_33;
  wire p_38_34;
  wire g_38_34;
  wire p_38_35;
  wire g_38_35;
  wire p_38_36;
  wire g_38_36;
  wire p_38_37;
  wire g_38_37;
  wire p_39_39;
  wire g_39_39;
 assign p_39_39 = a[39] ^ b[39];
 assign g_39_39 = a[39] & b[39];
  wire p_39_0;
  wire g_39_0;
  wire p_39_1;
  wire g_39_1;
  wire p_39_2;
  wire g_39_2;
  wire p_39_3;
  wire g_39_3;
  wire p_39_4;
  wire g_39_4;
  wire p_39_5;
  wire g_39_5;
  wire p_39_6;
  wire g_39_6;
  wire p_39_7;
  wire g_39_7;
  wire p_39_8;
  wire g_39_8;
  wire p_39_9;
  wire g_39_9;
  wire p_39_10;
  wire g_39_10;
  wire p_39_11;
  wire g_39_11;
  wire p_39_12;
  wire g_39_12;
  wire p_39_13;
  wire g_39_13;
  wire p_39_14;
  wire g_39_14;
  wire p_39_15;
  wire g_39_15;
  wire p_39_16;
  wire g_39_16;
  wire p_39_17;
  wire g_39_17;
  wire p_39_18;
  wire g_39_18;
  wire p_39_19;
  wire g_39_19;
  wire p_39_20;
  wire g_39_20;
  wire p_39_21;
  wire g_39_21;
  wire p_39_22;
  wire g_39_22;
  wire p_39_23;
  wire g_39_23;
  wire p_39_24;
  wire g_39_24;
  wire p_39_25;
  wire g_39_25;
  wire p_39_26;
  wire g_39_26;
  wire p_39_27;
  wire g_39_27;
  wire p_39_28;
  wire g_39_28;
  wire p_39_29;
  wire g_39_29;
  wire p_39_30;
  wire g_39_30;
  wire p_39_31;
  wire g_39_31;
  wire p_39_32;
  wire g_39_32;
  wire p_39_33;
  wire g_39_33;
  wire p_39_34;
  wire g_39_34;
  wire p_39_35;
  wire g_39_35;
  wire p_39_36;
  wire g_39_36;
  wire p_39_37;
  wire g_39_37;
  wire p_39_38;
  wire g_39_38;
  wire p_40_40;
  wire g_40_40;
 assign p_40_40 = a[40] ^ b[40];
 assign g_40_40 = a[40] & b[40];
  wire p_40_0;
  wire g_40_0;
  wire p_40_1;
  wire g_40_1;
  wire p_40_2;
  wire g_40_2;
  wire p_40_3;
  wire g_40_3;
  wire p_40_4;
  wire g_40_4;
  wire p_40_5;
  wire g_40_5;
  wire p_40_6;
  wire g_40_6;
  wire p_40_7;
  wire g_40_7;
  wire p_40_8;
  wire g_40_8;
  wire p_40_9;
  wire g_40_9;
  wire p_40_10;
  wire g_40_10;
  wire p_40_11;
  wire g_40_11;
  wire p_40_12;
  wire g_40_12;
  wire p_40_13;
  wire g_40_13;
  wire p_40_14;
  wire g_40_14;
  wire p_40_15;
  wire g_40_15;
  wire p_40_16;
  wire g_40_16;
  wire p_40_17;
  wire g_40_17;
  wire p_40_18;
  wire g_40_18;
  wire p_40_19;
  wire g_40_19;
  wire p_40_20;
  wire g_40_20;
  wire p_40_21;
  wire g_40_21;
  wire p_40_22;
  wire g_40_22;
  wire p_40_23;
  wire g_40_23;
  wire p_40_24;
  wire g_40_24;
  wire p_40_25;
  wire g_40_25;
  wire p_40_26;
  wire g_40_26;
  wire p_40_27;
  wire g_40_27;
  wire p_40_28;
  wire g_40_28;
  wire p_40_29;
  wire g_40_29;
  wire p_40_30;
  wire g_40_30;
  wire p_40_31;
  wire g_40_31;
  wire p_40_32;
  wire g_40_32;
  wire p_40_33;
  wire g_40_33;
  wire p_40_34;
  wire g_40_34;
  wire p_40_35;
  wire g_40_35;
  wire p_40_36;
  wire g_40_36;
  wire p_40_37;
  wire g_40_37;
  wire p_40_38;
  wire g_40_38;
  wire p_40_39;
  wire g_40_39;
  wire p_41_41;
  wire g_41_41;
 assign p_41_41 = a[41] ^ b[41];
 assign g_41_41 = a[41] & b[41];
  wire p_41_0;
  wire g_41_0;
  wire p_41_1;
  wire g_41_1;
  wire p_41_2;
  wire g_41_2;
  wire p_41_3;
  wire g_41_3;
  wire p_41_4;
  wire g_41_4;
  wire p_41_5;
  wire g_41_5;
  wire p_41_6;
  wire g_41_6;
  wire p_41_7;
  wire g_41_7;
  wire p_41_8;
  wire g_41_8;
  wire p_41_9;
  wire g_41_9;
  wire p_41_10;
  wire g_41_10;
  wire p_41_11;
  wire g_41_11;
  wire p_41_12;
  wire g_41_12;
  wire p_41_13;
  wire g_41_13;
  wire p_41_14;
  wire g_41_14;
  wire p_41_15;
  wire g_41_15;
  wire p_41_16;
  wire g_41_16;
  wire p_41_17;
  wire g_41_17;
  wire p_41_18;
  wire g_41_18;
  wire p_41_19;
  wire g_41_19;
  wire p_41_20;
  wire g_41_20;
  wire p_41_21;
  wire g_41_21;
  wire p_41_22;
  wire g_41_22;
  wire p_41_23;
  wire g_41_23;
  wire p_41_24;
  wire g_41_24;
  wire p_41_25;
  wire g_41_25;
  wire p_41_26;
  wire g_41_26;
  wire p_41_27;
  wire g_41_27;
  wire p_41_28;
  wire g_41_28;
  wire p_41_29;
  wire g_41_29;
  wire p_41_30;
  wire g_41_30;
  wire p_41_31;
  wire g_41_31;
  wire p_41_32;
  wire g_41_32;
  wire p_41_33;
  wire g_41_33;
  wire p_41_34;
  wire g_41_34;
  wire p_41_35;
  wire g_41_35;
  wire p_41_36;
  wire g_41_36;
  wire p_41_37;
  wire g_41_37;
  wire p_41_38;
  wire g_41_38;
  wire p_41_39;
  wire g_41_39;
  wire p_41_40;
  wire g_41_40;
  wire p_42_42;
  wire g_42_42;
 assign p_42_42 = a[42] ^ b[42];
 assign g_42_42 = a[42] & b[42];
  wire p_42_0;
  wire g_42_0;
  wire p_42_1;
  wire g_42_1;
  wire p_42_2;
  wire g_42_2;
  wire p_42_3;
  wire g_42_3;
  wire p_42_4;
  wire g_42_4;
  wire p_42_5;
  wire g_42_5;
  wire p_42_6;
  wire g_42_6;
  wire p_42_7;
  wire g_42_7;
  wire p_42_8;
  wire g_42_8;
  wire p_42_9;
  wire g_42_9;
  wire p_42_10;
  wire g_42_10;
  wire p_42_11;
  wire g_42_11;
  wire p_42_12;
  wire g_42_12;
  wire p_42_13;
  wire g_42_13;
  wire p_42_14;
  wire g_42_14;
  wire p_42_15;
  wire g_42_15;
  wire p_42_16;
  wire g_42_16;
  wire p_42_17;
  wire g_42_17;
  wire p_42_18;
  wire g_42_18;
  wire p_42_19;
  wire g_42_19;
  wire p_42_20;
  wire g_42_20;
  wire p_42_21;
  wire g_42_21;
  wire p_42_22;
  wire g_42_22;
  wire p_42_23;
  wire g_42_23;
  wire p_42_24;
  wire g_42_24;
  wire p_42_25;
  wire g_42_25;
  wire p_42_26;
  wire g_42_26;
  wire p_42_27;
  wire g_42_27;
  wire p_42_28;
  wire g_42_28;
  wire p_42_29;
  wire g_42_29;
  wire p_42_30;
  wire g_42_30;
  wire p_42_31;
  wire g_42_31;
  wire p_42_32;
  wire g_42_32;
  wire p_42_33;
  wire g_42_33;
  wire p_42_34;
  wire g_42_34;
  wire p_42_35;
  wire g_42_35;
  wire p_42_36;
  wire g_42_36;
  wire p_42_37;
  wire g_42_37;
  wire p_42_38;
  wire g_42_38;
  wire p_42_39;
  wire g_42_39;
  wire p_42_40;
  wire g_42_40;
  wire p_42_41;
  wire g_42_41;
  wire p_43_43;
  wire g_43_43;
 assign p_43_43 = a[43] ^ b[43];
 assign g_43_43 = a[43] & b[43];
  wire p_43_0;
  wire g_43_0;
  wire p_43_1;
  wire g_43_1;
  wire p_43_2;
  wire g_43_2;
  wire p_43_3;
  wire g_43_3;
  wire p_43_4;
  wire g_43_4;
  wire p_43_5;
  wire g_43_5;
  wire p_43_6;
  wire g_43_6;
  wire p_43_7;
  wire g_43_7;
  wire p_43_8;
  wire g_43_8;
  wire p_43_9;
  wire g_43_9;
  wire p_43_10;
  wire g_43_10;
  wire p_43_11;
  wire g_43_11;
  wire p_43_12;
  wire g_43_12;
  wire p_43_13;
  wire g_43_13;
  wire p_43_14;
  wire g_43_14;
  wire p_43_15;
  wire g_43_15;
  wire p_43_16;
  wire g_43_16;
  wire p_43_17;
  wire g_43_17;
  wire p_43_18;
  wire g_43_18;
  wire p_43_19;
  wire g_43_19;
  wire p_43_20;
  wire g_43_20;
  wire p_43_21;
  wire g_43_21;
  wire p_43_22;
  wire g_43_22;
  wire p_43_23;
  wire g_43_23;
  wire p_43_24;
  wire g_43_24;
  wire p_43_25;
  wire g_43_25;
  wire p_43_26;
  wire g_43_26;
  wire p_43_27;
  wire g_43_27;
  wire p_43_28;
  wire g_43_28;
  wire p_43_29;
  wire g_43_29;
  wire p_43_30;
  wire g_43_30;
  wire p_43_31;
  wire g_43_31;
  wire p_43_32;
  wire g_43_32;
  wire p_43_33;
  wire g_43_33;
  wire p_43_34;
  wire g_43_34;
  wire p_43_35;
  wire g_43_35;
  wire p_43_36;
  wire g_43_36;
  wire p_43_37;
  wire g_43_37;
  wire p_43_38;
  wire g_43_38;
  wire p_43_39;
  wire g_43_39;
  wire p_43_40;
  wire g_43_40;
  wire p_43_41;
  wire g_43_41;
  wire p_43_42;
  wire g_43_42;
  wire p_44_44;
  wire g_44_44;
 assign p_44_44 = a[44] ^ b[44];
 assign g_44_44 = a[44] & b[44];
  wire p_44_0;
  wire g_44_0;
  wire p_44_1;
  wire g_44_1;
  wire p_44_2;
  wire g_44_2;
  wire p_44_3;
  wire g_44_3;
  wire p_44_4;
  wire g_44_4;
  wire p_44_5;
  wire g_44_5;
  wire p_44_6;
  wire g_44_6;
  wire p_44_7;
  wire g_44_7;
  wire p_44_8;
  wire g_44_8;
  wire p_44_9;
  wire g_44_9;
  wire p_44_10;
  wire g_44_10;
  wire p_44_11;
  wire g_44_11;
  wire p_44_12;
  wire g_44_12;
  wire p_44_13;
  wire g_44_13;
  wire p_44_14;
  wire g_44_14;
  wire p_44_15;
  wire g_44_15;
  wire p_44_16;
  wire g_44_16;
  wire p_44_17;
  wire g_44_17;
  wire p_44_18;
  wire g_44_18;
  wire p_44_19;
  wire g_44_19;
  wire p_44_20;
  wire g_44_20;
  wire p_44_21;
  wire g_44_21;
  wire p_44_22;
  wire g_44_22;
  wire p_44_23;
  wire g_44_23;
  wire p_44_24;
  wire g_44_24;
  wire p_44_25;
  wire g_44_25;
  wire p_44_26;
  wire g_44_26;
  wire p_44_27;
  wire g_44_27;
  wire p_44_28;
  wire g_44_28;
  wire p_44_29;
  wire g_44_29;
  wire p_44_30;
  wire g_44_30;
  wire p_44_31;
  wire g_44_31;
  wire p_44_32;
  wire g_44_32;
  wire p_44_33;
  wire g_44_33;
  wire p_44_34;
  wire g_44_34;
  wire p_44_35;
  wire g_44_35;
  wire p_44_36;
  wire g_44_36;
  wire p_44_37;
  wire g_44_37;
  wire p_44_38;
  wire g_44_38;
  wire p_44_39;
  wire g_44_39;
  wire p_44_40;
  wire g_44_40;
  wire p_44_41;
  wire g_44_41;
  wire p_44_42;
  wire g_44_42;
  wire p_44_43;
  wire g_44_43;
  wire p_45_45;
  wire g_45_45;
 assign p_45_45 = a[45] ^ b[45];
 assign g_45_45 = a[45] & b[45];
  wire p_45_0;
  wire g_45_0;
  wire p_45_1;
  wire g_45_1;
  wire p_45_2;
  wire g_45_2;
  wire p_45_3;
  wire g_45_3;
  wire p_45_4;
  wire g_45_4;
  wire p_45_5;
  wire g_45_5;
  wire p_45_6;
  wire g_45_6;
  wire p_45_7;
  wire g_45_7;
  wire p_45_8;
  wire g_45_8;
  wire p_45_9;
  wire g_45_9;
  wire p_45_10;
  wire g_45_10;
  wire p_45_11;
  wire g_45_11;
  wire p_45_12;
  wire g_45_12;
  wire p_45_13;
  wire g_45_13;
  wire p_45_14;
  wire g_45_14;
  wire p_45_15;
  wire g_45_15;
  wire p_45_16;
  wire g_45_16;
  wire p_45_17;
  wire g_45_17;
  wire p_45_18;
  wire g_45_18;
  wire p_45_19;
  wire g_45_19;
  wire p_45_20;
  wire g_45_20;
  wire p_45_21;
  wire g_45_21;
  wire p_45_22;
  wire g_45_22;
  wire p_45_23;
  wire g_45_23;
  wire p_45_24;
  wire g_45_24;
  wire p_45_25;
  wire g_45_25;
  wire p_45_26;
  wire g_45_26;
  wire p_45_27;
  wire g_45_27;
  wire p_45_28;
  wire g_45_28;
  wire p_45_29;
  wire g_45_29;
  wire p_45_30;
  wire g_45_30;
  wire p_45_31;
  wire g_45_31;
  wire p_45_32;
  wire g_45_32;
  wire p_45_33;
  wire g_45_33;
  wire p_45_34;
  wire g_45_34;
  wire p_45_35;
  wire g_45_35;
  wire p_45_36;
  wire g_45_36;
  wire p_45_37;
  wire g_45_37;
  wire p_45_38;
  wire g_45_38;
  wire p_45_39;
  wire g_45_39;
  wire p_45_40;
  wire g_45_40;
  wire p_45_41;
  wire g_45_41;
  wire p_45_42;
  wire g_45_42;
  wire p_45_43;
  wire g_45_43;
  wire p_45_44;
  wire g_45_44;
  wire p_46_46;
  wire g_46_46;
 assign p_46_46 = a[46] ^ b[46];
 assign g_46_46 = a[46] & b[46];
  wire p_46_0;
  wire g_46_0;
  wire p_46_1;
  wire g_46_1;
  wire p_46_2;
  wire g_46_2;
  wire p_46_3;
  wire g_46_3;
  wire p_46_4;
  wire g_46_4;
  wire p_46_5;
  wire g_46_5;
  wire p_46_6;
  wire g_46_6;
  wire p_46_7;
  wire g_46_7;
  wire p_46_8;
  wire g_46_8;
  wire p_46_9;
  wire g_46_9;
  wire p_46_10;
  wire g_46_10;
  wire p_46_11;
  wire g_46_11;
  wire p_46_12;
  wire g_46_12;
  wire p_46_13;
  wire g_46_13;
  wire p_46_14;
  wire g_46_14;
  wire p_46_15;
  wire g_46_15;
  wire p_46_16;
  wire g_46_16;
  wire p_46_17;
  wire g_46_17;
  wire p_46_18;
  wire g_46_18;
  wire p_46_19;
  wire g_46_19;
  wire p_46_20;
  wire g_46_20;
  wire p_46_21;
  wire g_46_21;
  wire p_46_22;
  wire g_46_22;
  wire p_46_23;
  wire g_46_23;
  wire p_46_24;
  wire g_46_24;
  wire p_46_25;
  wire g_46_25;
  wire p_46_26;
  wire g_46_26;
  wire p_46_27;
  wire g_46_27;
  wire p_46_28;
  wire g_46_28;
  wire p_46_29;
  wire g_46_29;
  wire p_46_30;
  wire g_46_30;
  wire p_46_31;
  wire g_46_31;
  wire p_46_32;
  wire g_46_32;
  wire p_46_33;
  wire g_46_33;
  wire p_46_34;
  wire g_46_34;
  wire p_46_35;
  wire g_46_35;
  wire p_46_36;
  wire g_46_36;
  wire p_46_37;
  wire g_46_37;
  wire p_46_38;
  wire g_46_38;
  wire p_46_39;
  wire g_46_39;
  wire p_46_40;
  wire g_46_40;
  wire p_46_41;
  wire g_46_41;
  wire p_46_42;
  wire g_46_42;
  wire p_46_43;
  wire g_46_43;
  wire p_46_44;
  wire g_46_44;
  wire p_46_45;
  wire g_46_45;
  wire p_47_47;
  wire g_47_47;
 assign p_47_47 = a[47] ^ b[47];
 assign g_47_47 = a[47] & b[47];
  wire p_47_0;
  wire g_47_0;
  wire p_47_1;
  wire g_47_1;
  wire p_47_2;
  wire g_47_2;
  wire p_47_3;
  wire g_47_3;
  wire p_47_4;
  wire g_47_4;
  wire p_47_5;
  wire g_47_5;
  wire p_47_6;
  wire g_47_6;
  wire p_47_7;
  wire g_47_7;
  wire p_47_8;
  wire g_47_8;
  wire p_47_9;
  wire g_47_9;
  wire p_47_10;
  wire g_47_10;
  wire p_47_11;
  wire g_47_11;
  wire p_47_12;
  wire g_47_12;
  wire p_47_13;
  wire g_47_13;
  wire p_47_14;
  wire g_47_14;
  wire p_47_15;
  wire g_47_15;
  wire p_47_16;
  wire g_47_16;
  wire p_47_17;
  wire g_47_17;
  wire p_47_18;
  wire g_47_18;
  wire p_47_19;
  wire g_47_19;
  wire p_47_20;
  wire g_47_20;
  wire p_47_21;
  wire g_47_21;
  wire p_47_22;
  wire g_47_22;
  wire p_47_23;
  wire g_47_23;
  wire p_47_24;
  wire g_47_24;
  wire p_47_25;
  wire g_47_25;
  wire p_47_26;
  wire g_47_26;
  wire p_47_27;
  wire g_47_27;
  wire p_47_28;
  wire g_47_28;
  wire p_47_29;
  wire g_47_29;
  wire p_47_30;
  wire g_47_30;
  wire p_47_31;
  wire g_47_31;
  wire p_47_32;
  wire g_47_32;
  wire p_47_33;
  wire g_47_33;
  wire p_47_34;
  wire g_47_34;
  wire p_47_35;
  wire g_47_35;
  wire p_47_36;
  wire g_47_36;
  wire p_47_37;
  wire g_47_37;
  wire p_47_38;
  wire g_47_38;
  wire p_47_39;
  wire g_47_39;
  wire p_47_40;
  wire g_47_40;
  wire p_47_41;
  wire g_47_41;
  wire p_47_42;
  wire g_47_42;
  wire p_47_43;
  wire g_47_43;
  wire p_47_44;
  wire g_47_44;
  wire p_47_45;
  wire g_47_45;
  wire p_47_46;
  wire g_47_46;
  wire p_48_48;
  wire g_48_48;
 assign p_48_48 = a[48] ^ b[48];
 assign g_48_48 = a[48] & b[48];
  wire p_48_0;
  wire g_48_0;
  wire p_48_1;
  wire g_48_1;
  wire p_48_2;
  wire g_48_2;
  wire p_48_3;
  wire g_48_3;
  wire p_48_4;
  wire g_48_4;
  wire p_48_5;
  wire g_48_5;
  wire p_48_6;
  wire g_48_6;
  wire p_48_7;
  wire g_48_7;
  wire p_48_8;
  wire g_48_8;
  wire p_48_9;
  wire g_48_9;
  wire p_48_10;
  wire g_48_10;
  wire p_48_11;
  wire g_48_11;
  wire p_48_12;
  wire g_48_12;
  wire p_48_13;
  wire g_48_13;
  wire p_48_14;
  wire g_48_14;
  wire p_48_15;
  wire g_48_15;
  wire p_48_16;
  wire g_48_16;
  wire p_48_17;
  wire g_48_17;
  wire p_48_18;
  wire g_48_18;
  wire p_48_19;
  wire g_48_19;
  wire p_48_20;
  wire g_48_20;
  wire p_48_21;
  wire g_48_21;
  wire p_48_22;
  wire g_48_22;
  wire p_48_23;
  wire g_48_23;
  wire p_48_24;
  wire g_48_24;
  wire p_48_25;
  wire g_48_25;
  wire p_48_26;
  wire g_48_26;
  wire p_48_27;
  wire g_48_27;
  wire p_48_28;
  wire g_48_28;
  wire p_48_29;
  wire g_48_29;
  wire p_48_30;
  wire g_48_30;
  wire p_48_31;
  wire g_48_31;
  wire p_48_32;
  wire g_48_32;
  wire p_48_33;
  wire g_48_33;
  wire p_48_34;
  wire g_48_34;
  wire p_48_35;
  wire g_48_35;
  wire p_48_36;
  wire g_48_36;
  wire p_48_37;
  wire g_48_37;
  wire p_48_38;
  wire g_48_38;
  wire p_48_39;
  wire g_48_39;
  wire p_48_40;
  wire g_48_40;
  wire p_48_41;
  wire g_48_41;
  wire p_48_42;
  wire g_48_42;
  wire p_48_43;
  wire g_48_43;
  wire p_48_44;
  wire g_48_44;
  wire p_48_45;
  wire g_48_45;
  wire p_48_46;
  wire g_48_46;
  wire p_48_47;
  wire g_48_47;
  wire p_49_49;
  wire g_49_49;
 assign p_49_49 = a[49] ^ b[49];
 assign g_49_49 = a[49] & b[49];
  wire p_49_0;
  wire g_49_0;
  wire p_49_1;
  wire g_49_1;
  wire p_49_2;
  wire g_49_2;
  wire p_49_3;
  wire g_49_3;
  wire p_49_4;
  wire g_49_4;
  wire p_49_5;
  wire g_49_5;
  wire p_49_6;
  wire g_49_6;
  wire p_49_7;
  wire g_49_7;
  wire p_49_8;
  wire g_49_8;
  wire p_49_9;
  wire g_49_9;
  wire p_49_10;
  wire g_49_10;
  wire p_49_11;
  wire g_49_11;
  wire p_49_12;
  wire g_49_12;
  wire p_49_13;
  wire g_49_13;
  wire p_49_14;
  wire g_49_14;
  wire p_49_15;
  wire g_49_15;
  wire p_49_16;
  wire g_49_16;
  wire p_49_17;
  wire g_49_17;
  wire p_49_18;
  wire g_49_18;
  wire p_49_19;
  wire g_49_19;
  wire p_49_20;
  wire g_49_20;
  wire p_49_21;
  wire g_49_21;
  wire p_49_22;
  wire g_49_22;
  wire p_49_23;
  wire g_49_23;
  wire p_49_24;
  wire g_49_24;
  wire p_49_25;
  wire g_49_25;
  wire p_49_26;
  wire g_49_26;
  wire p_49_27;
  wire g_49_27;
  wire p_49_28;
  wire g_49_28;
  wire p_49_29;
  wire g_49_29;
  wire p_49_30;
  wire g_49_30;
  wire p_49_31;
  wire g_49_31;
  wire p_49_32;
  wire g_49_32;
  wire p_49_33;
  wire g_49_33;
  wire p_49_34;
  wire g_49_34;
  wire p_49_35;
  wire g_49_35;
  wire p_49_36;
  wire g_49_36;
  wire p_49_37;
  wire g_49_37;
  wire p_49_38;
  wire g_49_38;
  wire p_49_39;
  wire g_49_39;
  wire p_49_40;
  wire g_49_40;
  wire p_49_41;
  wire g_49_41;
  wire p_49_42;
  wire g_49_42;
  wire p_49_43;
  wire g_49_43;
  wire p_49_44;
  wire g_49_44;
  wire p_49_45;
  wire g_49_45;
  wire p_49_46;
  wire g_49_46;
  wire p_49_47;
  wire g_49_47;
  wire p_49_48;
  wire g_49_48;
  wire p_50_50;
  wire g_50_50;
 assign p_50_50 = a[50] ^ b[50];
 assign g_50_50 = a[50] & b[50];
  wire p_50_0;
  wire g_50_0;
  wire p_50_1;
  wire g_50_1;
  wire p_50_2;
  wire g_50_2;
  wire p_50_3;
  wire g_50_3;
  wire p_50_4;
  wire g_50_4;
  wire p_50_5;
  wire g_50_5;
  wire p_50_6;
  wire g_50_6;
  wire p_50_7;
  wire g_50_7;
  wire p_50_8;
  wire g_50_8;
  wire p_50_9;
  wire g_50_9;
  wire p_50_10;
  wire g_50_10;
  wire p_50_11;
  wire g_50_11;
  wire p_50_12;
  wire g_50_12;
  wire p_50_13;
  wire g_50_13;
  wire p_50_14;
  wire g_50_14;
  wire p_50_15;
  wire g_50_15;
  wire p_50_16;
  wire g_50_16;
  wire p_50_17;
  wire g_50_17;
  wire p_50_18;
  wire g_50_18;
  wire p_50_19;
  wire g_50_19;
  wire p_50_20;
  wire g_50_20;
  wire p_50_21;
  wire g_50_21;
  wire p_50_22;
  wire g_50_22;
  wire p_50_23;
  wire g_50_23;
  wire p_50_24;
  wire g_50_24;
  wire p_50_25;
  wire g_50_25;
  wire p_50_26;
  wire g_50_26;
  wire p_50_27;
  wire g_50_27;
  wire p_50_28;
  wire g_50_28;
  wire p_50_29;
  wire g_50_29;
  wire p_50_30;
  wire g_50_30;
  wire p_50_31;
  wire g_50_31;
  wire p_50_32;
  wire g_50_32;
  wire p_50_33;
  wire g_50_33;
  wire p_50_34;
  wire g_50_34;
  wire p_50_35;
  wire g_50_35;
  wire p_50_36;
  wire g_50_36;
  wire p_50_37;
  wire g_50_37;
  wire p_50_38;
  wire g_50_38;
  wire p_50_39;
  wire g_50_39;
  wire p_50_40;
  wire g_50_40;
  wire p_50_41;
  wire g_50_41;
  wire p_50_42;
  wire g_50_42;
  wire p_50_43;
  wire g_50_43;
  wire p_50_44;
  wire g_50_44;
  wire p_50_45;
  wire g_50_45;
  wire p_50_46;
  wire g_50_46;
  wire p_50_47;
  wire g_50_47;
  wire p_50_48;
  wire g_50_48;
  wire p_50_49;
  wire g_50_49;
  wire p_51_51;
  wire g_51_51;
 assign p_51_51 = a[51] ^ b[51];
 assign g_51_51 = a[51] & b[51];
  wire p_51_0;
  wire g_51_0;
  wire p_51_1;
  wire g_51_1;
  wire p_51_2;
  wire g_51_2;
  wire p_51_3;
  wire g_51_3;
  wire p_51_4;
  wire g_51_4;
  wire p_51_5;
  wire g_51_5;
  wire p_51_6;
  wire g_51_6;
  wire p_51_7;
  wire g_51_7;
  wire p_51_8;
  wire g_51_8;
  wire p_51_9;
  wire g_51_9;
  wire p_51_10;
  wire g_51_10;
  wire p_51_11;
  wire g_51_11;
  wire p_51_12;
  wire g_51_12;
  wire p_51_13;
  wire g_51_13;
  wire p_51_14;
  wire g_51_14;
  wire p_51_15;
  wire g_51_15;
  wire p_51_16;
  wire g_51_16;
  wire p_51_17;
  wire g_51_17;
  wire p_51_18;
  wire g_51_18;
  wire p_51_19;
  wire g_51_19;
  wire p_51_20;
  wire g_51_20;
  wire p_51_21;
  wire g_51_21;
  wire p_51_22;
  wire g_51_22;
  wire p_51_23;
  wire g_51_23;
  wire p_51_24;
  wire g_51_24;
  wire p_51_25;
  wire g_51_25;
  wire p_51_26;
  wire g_51_26;
  wire p_51_27;
  wire g_51_27;
  wire p_51_28;
  wire g_51_28;
  wire p_51_29;
  wire g_51_29;
  wire p_51_30;
  wire g_51_30;
  wire p_51_31;
  wire g_51_31;
  wire p_51_32;
  wire g_51_32;
  wire p_51_33;
  wire g_51_33;
  wire p_51_34;
  wire g_51_34;
  wire p_51_35;
  wire g_51_35;
  wire p_51_36;
  wire g_51_36;
  wire p_51_37;
  wire g_51_37;
  wire p_51_38;
  wire g_51_38;
  wire p_51_39;
  wire g_51_39;
  wire p_51_40;
  wire g_51_40;
  wire p_51_41;
  wire g_51_41;
  wire p_51_42;
  wire g_51_42;
  wire p_51_43;
  wire g_51_43;
  wire p_51_44;
  wire g_51_44;
  wire p_51_45;
  wire g_51_45;
  wire p_51_46;
  wire g_51_46;
  wire p_51_47;
  wire g_51_47;
  wire p_51_48;
  wire g_51_48;
  wire p_51_49;
  wire g_51_49;
  wire p_51_50;
  wire g_51_50;
  wire p_52_52;
  wire g_52_52;
 assign p_52_52 = a[52] ^ b[52];
 assign g_52_52 = a[52] & b[52];
  wire p_52_0;
  wire g_52_0;
  wire p_52_1;
  wire g_52_1;
  wire p_52_2;
  wire g_52_2;
  wire p_52_3;
  wire g_52_3;
  wire p_52_4;
  wire g_52_4;
  wire p_52_5;
  wire g_52_5;
  wire p_52_6;
  wire g_52_6;
  wire p_52_7;
  wire g_52_7;
  wire p_52_8;
  wire g_52_8;
  wire p_52_9;
  wire g_52_9;
  wire p_52_10;
  wire g_52_10;
  wire p_52_11;
  wire g_52_11;
  wire p_52_12;
  wire g_52_12;
  wire p_52_13;
  wire g_52_13;
  wire p_52_14;
  wire g_52_14;
  wire p_52_15;
  wire g_52_15;
  wire p_52_16;
  wire g_52_16;
  wire p_52_17;
  wire g_52_17;
  wire p_52_18;
  wire g_52_18;
  wire p_52_19;
  wire g_52_19;
  wire p_52_20;
  wire g_52_20;
  wire p_52_21;
  wire g_52_21;
  wire p_52_22;
  wire g_52_22;
  wire p_52_23;
  wire g_52_23;
  wire p_52_24;
  wire g_52_24;
  wire p_52_25;
  wire g_52_25;
  wire p_52_26;
  wire g_52_26;
  wire p_52_27;
  wire g_52_27;
  wire p_52_28;
  wire g_52_28;
  wire p_52_29;
  wire g_52_29;
  wire p_52_30;
  wire g_52_30;
  wire p_52_31;
  wire g_52_31;
  wire p_52_32;
  wire g_52_32;
  wire p_52_33;
  wire g_52_33;
  wire p_52_34;
  wire g_52_34;
  wire p_52_35;
  wire g_52_35;
  wire p_52_36;
  wire g_52_36;
  wire p_52_37;
  wire g_52_37;
  wire p_52_38;
  wire g_52_38;
  wire p_52_39;
  wire g_52_39;
  wire p_52_40;
  wire g_52_40;
  wire p_52_41;
  wire g_52_41;
  wire p_52_42;
  wire g_52_42;
  wire p_52_43;
  wire g_52_43;
  wire p_52_44;
  wire g_52_44;
  wire p_52_45;
  wire g_52_45;
  wire p_52_46;
  wire g_52_46;
  wire p_52_47;
  wire g_52_47;
  wire p_52_48;
  wire g_52_48;
  wire p_52_49;
  wire g_52_49;
  wire p_52_50;
  wire g_52_50;
  wire p_52_51;
  wire g_52_51;
  wire p_53_53;
  wire g_53_53;
 assign p_53_53 = a[53] ^ b[53];
 assign g_53_53 = a[53] & b[53];
  wire p_53_0;
  wire g_53_0;
  wire p_53_1;
  wire g_53_1;
  wire p_53_2;
  wire g_53_2;
  wire p_53_3;
  wire g_53_3;
  wire p_53_4;
  wire g_53_4;
  wire p_53_5;
  wire g_53_5;
  wire p_53_6;
  wire g_53_6;
  wire p_53_7;
  wire g_53_7;
  wire p_53_8;
  wire g_53_8;
  wire p_53_9;
  wire g_53_9;
  wire p_53_10;
  wire g_53_10;
  wire p_53_11;
  wire g_53_11;
  wire p_53_12;
  wire g_53_12;
  wire p_53_13;
  wire g_53_13;
  wire p_53_14;
  wire g_53_14;
  wire p_53_15;
  wire g_53_15;
  wire p_53_16;
  wire g_53_16;
  wire p_53_17;
  wire g_53_17;
  wire p_53_18;
  wire g_53_18;
  wire p_53_19;
  wire g_53_19;
  wire p_53_20;
  wire g_53_20;
  wire p_53_21;
  wire g_53_21;
  wire p_53_22;
  wire g_53_22;
  wire p_53_23;
  wire g_53_23;
  wire p_53_24;
  wire g_53_24;
  wire p_53_25;
  wire g_53_25;
  wire p_53_26;
  wire g_53_26;
  wire p_53_27;
  wire g_53_27;
  wire p_53_28;
  wire g_53_28;
  wire p_53_29;
  wire g_53_29;
  wire p_53_30;
  wire g_53_30;
  wire p_53_31;
  wire g_53_31;
  wire p_53_32;
  wire g_53_32;
  wire p_53_33;
  wire g_53_33;
  wire p_53_34;
  wire g_53_34;
  wire p_53_35;
  wire g_53_35;
  wire p_53_36;
  wire g_53_36;
  wire p_53_37;
  wire g_53_37;
  wire p_53_38;
  wire g_53_38;
  wire p_53_39;
  wire g_53_39;
  wire p_53_40;
  wire g_53_40;
  wire p_53_41;
  wire g_53_41;
  wire p_53_42;
  wire g_53_42;
  wire p_53_43;
  wire g_53_43;
  wire p_53_44;
  wire g_53_44;
  wire p_53_45;
  wire g_53_45;
  wire p_53_46;
  wire g_53_46;
  wire p_53_47;
  wire g_53_47;
  wire p_53_48;
  wire g_53_48;
  wire p_53_49;
  wire g_53_49;
  wire p_53_50;
  wire g_53_50;
  wire p_53_51;
  wire g_53_51;
  wire p_53_52;
  wire g_53_52;
  wire p_54_54;
  wire g_54_54;
 assign p_54_54 = a[54] ^ b[54];
 assign g_54_54 = a[54] & b[54];
  wire p_54_0;
  wire g_54_0;
  wire p_54_1;
  wire g_54_1;
  wire p_54_2;
  wire g_54_2;
  wire p_54_3;
  wire g_54_3;
  wire p_54_4;
  wire g_54_4;
  wire p_54_5;
  wire g_54_5;
  wire p_54_6;
  wire g_54_6;
  wire p_54_7;
  wire g_54_7;
  wire p_54_8;
  wire g_54_8;
  wire p_54_9;
  wire g_54_9;
  wire p_54_10;
  wire g_54_10;
  wire p_54_11;
  wire g_54_11;
  wire p_54_12;
  wire g_54_12;
  wire p_54_13;
  wire g_54_13;
  wire p_54_14;
  wire g_54_14;
  wire p_54_15;
  wire g_54_15;
  wire p_54_16;
  wire g_54_16;
  wire p_54_17;
  wire g_54_17;
  wire p_54_18;
  wire g_54_18;
  wire p_54_19;
  wire g_54_19;
  wire p_54_20;
  wire g_54_20;
  wire p_54_21;
  wire g_54_21;
  wire p_54_22;
  wire g_54_22;
  wire p_54_23;
  wire g_54_23;
  wire p_54_24;
  wire g_54_24;
  wire p_54_25;
  wire g_54_25;
  wire p_54_26;
  wire g_54_26;
  wire p_54_27;
  wire g_54_27;
  wire p_54_28;
  wire g_54_28;
  wire p_54_29;
  wire g_54_29;
  wire p_54_30;
  wire g_54_30;
  wire p_54_31;
  wire g_54_31;
  wire p_54_32;
  wire g_54_32;
  wire p_54_33;
  wire g_54_33;
  wire p_54_34;
  wire g_54_34;
  wire p_54_35;
  wire g_54_35;
  wire p_54_36;
  wire g_54_36;
  wire p_54_37;
  wire g_54_37;
  wire p_54_38;
  wire g_54_38;
  wire p_54_39;
  wire g_54_39;
  wire p_54_40;
  wire g_54_40;
  wire p_54_41;
  wire g_54_41;
  wire p_54_42;
  wire g_54_42;
  wire p_54_43;
  wire g_54_43;
  wire p_54_44;
  wire g_54_44;
  wire p_54_45;
  wire g_54_45;
  wire p_54_46;
  wire g_54_46;
  wire p_54_47;
  wire g_54_47;
  wire p_54_48;
  wire g_54_48;
  wire p_54_49;
  wire g_54_49;
  wire p_54_50;
  wire g_54_50;
  wire p_54_51;
  wire g_54_51;
  wire p_54_52;
  wire g_54_52;
  wire p_54_53;
  wire g_54_53;
  wire p_55_55;
  wire g_55_55;
 assign p_55_55 = a[55] ^ b[55];
 assign g_55_55 = a[55] & b[55];
  wire p_55_0;
  wire g_55_0;
  wire p_55_1;
  wire g_55_1;
  wire p_55_2;
  wire g_55_2;
  wire p_55_3;
  wire g_55_3;
  wire p_55_4;
  wire g_55_4;
  wire p_55_5;
  wire g_55_5;
  wire p_55_6;
  wire g_55_6;
  wire p_55_7;
  wire g_55_7;
  wire p_55_8;
  wire g_55_8;
  wire p_55_9;
  wire g_55_9;
  wire p_55_10;
  wire g_55_10;
  wire p_55_11;
  wire g_55_11;
  wire p_55_12;
  wire g_55_12;
  wire p_55_13;
  wire g_55_13;
  wire p_55_14;
  wire g_55_14;
  wire p_55_15;
  wire g_55_15;
  wire p_55_16;
  wire g_55_16;
  wire p_55_17;
  wire g_55_17;
  wire p_55_18;
  wire g_55_18;
  wire p_55_19;
  wire g_55_19;
  wire p_55_20;
  wire g_55_20;
  wire p_55_21;
  wire g_55_21;
  wire p_55_22;
  wire g_55_22;
  wire p_55_23;
  wire g_55_23;
  wire p_55_24;
  wire g_55_24;
  wire p_55_25;
  wire g_55_25;
  wire p_55_26;
  wire g_55_26;
  wire p_55_27;
  wire g_55_27;
  wire p_55_28;
  wire g_55_28;
  wire p_55_29;
  wire g_55_29;
  wire p_55_30;
  wire g_55_30;
  wire p_55_31;
  wire g_55_31;
  wire p_55_32;
  wire g_55_32;
  wire p_55_33;
  wire g_55_33;
  wire p_55_34;
  wire g_55_34;
  wire p_55_35;
  wire g_55_35;
  wire p_55_36;
  wire g_55_36;
  wire p_55_37;
  wire g_55_37;
  wire p_55_38;
  wire g_55_38;
  wire p_55_39;
  wire g_55_39;
  wire p_55_40;
  wire g_55_40;
  wire p_55_41;
  wire g_55_41;
  wire p_55_42;
  wire g_55_42;
  wire p_55_43;
  wire g_55_43;
  wire p_55_44;
  wire g_55_44;
  wire p_55_45;
  wire g_55_45;
  wire p_55_46;
  wire g_55_46;
  wire p_55_47;
  wire g_55_47;
  wire p_55_48;
  wire g_55_48;
  wire p_55_49;
  wire g_55_49;
  wire p_55_50;
  wire g_55_50;
  wire p_55_51;
  wire g_55_51;
  wire p_55_52;
  wire g_55_52;
  wire p_55_53;
  wire g_55_53;
  wire p_55_54;
  wire g_55_54;
  wire p_56_56;
  wire g_56_56;
 assign p_56_56 = a[56] ^ b[56];
 assign g_56_56 = a[56] & b[56];
  wire p_56_0;
  wire g_56_0;
  wire p_56_1;
  wire g_56_1;
  wire p_56_2;
  wire g_56_2;
  wire p_56_3;
  wire g_56_3;
  wire p_56_4;
  wire g_56_4;
  wire p_56_5;
  wire g_56_5;
  wire p_56_6;
  wire g_56_6;
  wire p_56_7;
  wire g_56_7;
  wire p_56_8;
  wire g_56_8;
  wire p_56_9;
  wire g_56_9;
  wire p_56_10;
  wire g_56_10;
  wire p_56_11;
  wire g_56_11;
  wire p_56_12;
  wire g_56_12;
  wire p_56_13;
  wire g_56_13;
  wire p_56_14;
  wire g_56_14;
  wire p_56_15;
  wire g_56_15;
  wire p_56_16;
  wire g_56_16;
  wire p_56_17;
  wire g_56_17;
  wire p_56_18;
  wire g_56_18;
  wire p_56_19;
  wire g_56_19;
  wire p_56_20;
  wire g_56_20;
  wire p_56_21;
  wire g_56_21;
  wire p_56_22;
  wire g_56_22;
  wire p_56_23;
  wire g_56_23;
  wire p_56_24;
  wire g_56_24;
  wire p_56_25;
  wire g_56_25;
  wire p_56_26;
  wire g_56_26;
  wire p_56_27;
  wire g_56_27;
  wire p_56_28;
  wire g_56_28;
  wire p_56_29;
  wire g_56_29;
  wire p_56_30;
  wire g_56_30;
  wire p_56_31;
  wire g_56_31;
  wire p_56_32;
  wire g_56_32;
  wire p_56_33;
  wire g_56_33;
  wire p_56_34;
  wire g_56_34;
  wire p_56_35;
  wire g_56_35;
  wire p_56_36;
  wire g_56_36;
  wire p_56_37;
  wire g_56_37;
  wire p_56_38;
  wire g_56_38;
  wire p_56_39;
  wire g_56_39;
  wire p_56_40;
  wire g_56_40;
  wire p_56_41;
  wire g_56_41;
  wire p_56_42;
  wire g_56_42;
  wire p_56_43;
  wire g_56_43;
  wire p_56_44;
  wire g_56_44;
  wire p_56_45;
  wire g_56_45;
  wire p_56_46;
  wire g_56_46;
  wire p_56_47;
  wire g_56_47;
  wire p_56_48;
  wire g_56_48;
  wire p_56_49;
  wire g_56_49;
  wire p_56_50;
  wire g_56_50;
  wire p_56_51;
  wire g_56_51;
  wire p_56_52;
  wire g_56_52;
  wire p_56_53;
  wire g_56_53;
  wire p_56_54;
  wire g_56_54;
  wire p_56_55;
  wire g_56_55;
  wire p_57_57;
  wire g_57_57;
 assign p_57_57 = a[57] ^ b[57];
 assign g_57_57 = a[57] & b[57];
  wire p_57_0;
  wire g_57_0;
  wire p_57_1;
  wire g_57_1;
  wire p_57_2;
  wire g_57_2;
  wire p_57_3;
  wire g_57_3;
  wire p_57_4;
  wire g_57_4;
  wire p_57_5;
  wire g_57_5;
  wire p_57_6;
  wire g_57_6;
  wire p_57_7;
  wire g_57_7;
  wire p_57_8;
  wire g_57_8;
  wire p_57_9;
  wire g_57_9;
  wire p_57_10;
  wire g_57_10;
  wire p_57_11;
  wire g_57_11;
  wire p_57_12;
  wire g_57_12;
  wire p_57_13;
  wire g_57_13;
  wire p_57_14;
  wire g_57_14;
  wire p_57_15;
  wire g_57_15;
  wire p_57_16;
  wire g_57_16;
  wire p_57_17;
  wire g_57_17;
  wire p_57_18;
  wire g_57_18;
  wire p_57_19;
  wire g_57_19;
  wire p_57_20;
  wire g_57_20;
  wire p_57_21;
  wire g_57_21;
  wire p_57_22;
  wire g_57_22;
  wire p_57_23;
  wire g_57_23;
  wire p_57_24;
  wire g_57_24;
  wire p_57_25;
  wire g_57_25;
  wire p_57_26;
  wire g_57_26;
  wire p_57_27;
  wire g_57_27;
  wire p_57_28;
  wire g_57_28;
  wire p_57_29;
  wire g_57_29;
  wire p_57_30;
  wire g_57_30;
  wire p_57_31;
  wire g_57_31;
  wire p_57_32;
  wire g_57_32;
  wire p_57_33;
  wire g_57_33;
  wire p_57_34;
  wire g_57_34;
  wire p_57_35;
  wire g_57_35;
  wire p_57_36;
  wire g_57_36;
  wire p_57_37;
  wire g_57_37;
  wire p_57_38;
  wire g_57_38;
  wire p_57_39;
  wire g_57_39;
  wire p_57_40;
  wire g_57_40;
  wire p_57_41;
  wire g_57_41;
  wire p_57_42;
  wire g_57_42;
  wire p_57_43;
  wire g_57_43;
  wire p_57_44;
  wire g_57_44;
  wire p_57_45;
  wire g_57_45;
  wire p_57_46;
  wire g_57_46;
  wire p_57_47;
  wire g_57_47;
  wire p_57_48;
  wire g_57_48;
  wire p_57_49;
  wire g_57_49;
  wire p_57_50;
  wire g_57_50;
  wire p_57_51;
  wire g_57_51;
  wire p_57_52;
  wire g_57_52;
  wire p_57_53;
  wire g_57_53;
  wire p_57_54;
  wire g_57_54;
  wire p_57_55;
  wire g_57_55;
  wire p_57_56;
  wire g_57_56;
  wire p_58_58;
  wire g_58_58;
 assign p_58_58 = a[58] ^ b[58];
 assign g_58_58 = a[58] & b[58];
  wire p_58_0;
  wire g_58_0;
  wire p_58_1;
  wire g_58_1;
  wire p_58_2;
  wire g_58_2;
  wire p_58_3;
  wire g_58_3;
  wire p_58_4;
  wire g_58_4;
  wire p_58_5;
  wire g_58_5;
  wire p_58_6;
  wire g_58_6;
  wire p_58_7;
  wire g_58_7;
  wire p_58_8;
  wire g_58_8;
  wire p_58_9;
  wire g_58_9;
  wire p_58_10;
  wire g_58_10;
  wire p_58_11;
  wire g_58_11;
  wire p_58_12;
  wire g_58_12;
  wire p_58_13;
  wire g_58_13;
  wire p_58_14;
  wire g_58_14;
  wire p_58_15;
  wire g_58_15;
  wire p_58_16;
  wire g_58_16;
  wire p_58_17;
  wire g_58_17;
  wire p_58_18;
  wire g_58_18;
  wire p_58_19;
  wire g_58_19;
  wire p_58_20;
  wire g_58_20;
  wire p_58_21;
  wire g_58_21;
  wire p_58_22;
  wire g_58_22;
  wire p_58_23;
  wire g_58_23;
  wire p_58_24;
  wire g_58_24;
  wire p_58_25;
  wire g_58_25;
  wire p_58_26;
  wire g_58_26;
  wire p_58_27;
  wire g_58_27;
  wire p_58_28;
  wire g_58_28;
  wire p_58_29;
  wire g_58_29;
  wire p_58_30;
  wire g_58_30;
  wire p_58_31;
  wire g_58_31;
  wire p_58_32;
  wire g_58_32;
  wire p_58_33;
  wire g_58_33;
  wire p_58_34;
  wire g_58_34;
  wire p_58_35;
  wire g_58_35;
  wire p_58_36;
  wire g_58_36;
  wire p_58_37;
  wire g_58_37;
  wire p_58_38;
  wire g_58_38;
  wire p_58_39;
  wire g_58_39;
  wire p_58_40;
  wire g_58_40;
  wire p_58_41;
  wire g_58_41;
  wire p_58_42;
  wire g_58_42;
  wire p_58_43;
  wire g_58_43;
  wire p_58_44;
  wire g_58_44;
  wire p_58_45;
  wire g_58_45;
  wire p_58_46;
  wire g_58_46;
  wire p_58_47;
  wire g_58_47;
  wire p_58_48;
  wire g_58_48;
  wire p_58_49;
  wire g_58_49;
  wire p_58_50;
  wire g_58_50;
  wire p_58_51;
  wire g_58_51;
  wire p_58_52;
  wire g_58_52;
  wire p_58_53;
  wire g_58_53;
  wire p_58_54;
  wire g_58_54;
  wire p_58_55;
  wire g_58_55;
  wire p_58_56;
  wire g_58_56;
  wire p_58_57;
  wire g_58_57;
  wire p_59_59;
  wire g_59_59;
 assign p_59_59 = a[59] ^ b[59];
 assign g_59_59 = a[59] & b[59];
  wire p_59_0;
  wire g_59_0;
  wire p_59_1;
  wire g_59_1;
  wire p_59_2;
  wire g_59_2;
  wire p_59_3;
  wire g_59_3;
  wire p_59_4;
  wire g_59_4;
  wire p_59_5;
  wire g_59_5;
  wire p_59_6;
  wire g_59_6;
  wire p_59_7;
  wire g_59_7;
  wire p_59_8;
  wire g_59_8;
  wire p_59_9;
  wire g_59_9;
  wire p_59_10;
  wire g_59_10;
  wire p_59_11;
  wire g_59_11;
  wire p_59_12;
  wire g_59_12;
  wire p_59_13;
  wire g_59_13;
  wire p_59_14;
  wire g_59_14;
  wire p_59_15;
  wire g_59_15;
  wire p_59_16;
  wire g_59_16;
  wire p_59_17;
  wire g_59_17;
  wire p_59_18;
  wire g_59_18;
  wire p_59_19;
  wire g_59_19;
  wire p_59_20;
  wire g_59_20;
  wire p_59_21;
  wire g_59_21;
  wire p_59_22;
  wire g_59_22;
  wire p_59_23;
  wire g_59_23;
  wire p_59_24;
  wire g_59_24;
  wire p_59_25;
  wire g_59_25;
  wire p_59_26;
  wire g_59_26;
  wire p_59_27;
  wire g_59_27;
  wire p_59_28;
  wire g_59_28;
  wire p_59_29;
  wire g_59_29;
  wire p_59_30;
  wire g_59_30;
  wire p_59_31;
  wire g_59_31;
  wire p_59_32;
  wire g_59_32;
  wire p_59_33;
  wire g_59_33;
  wire p_59_34;
  wire g_59_34;
  wire p_59_35;
  wire g_59_35;
  wire p_59_36;
  wire g_59_36;
  wire p_59_37;
  wire g_59_37;
  wire p_59_38;
  wire g_59_38;
  wire p_59_39;
  wire g_59_39;
  wire p_59_40;
  wire g_59_40;
  wire p_59_41;
  wire g_59_41;
  wire p_59_42;
  wire g_59_42;
  wire p_59_43;
  wire g_59_43;
  wire p_59_44;
  wire g_59_44;
  wire p_59_45;
  wire g_59_45;
  wire p_59_46;
  wire g_59_46;
  wire p_59_47;
  wire g_59_47;
  wire p_59_48;
  wire g_59_48;
  wire p_59_49;
  wire g_59_49;
  wire p_59_50;
  wire g_59_50;
  wire p_59_51;
  wire g_59_51;
  wire p_59_52;
  wire g_59_52;
  wire p_59_53;
  wire g_59_53;
  wire p_59_54;
  wire g_59_54;
  wire p_59_55;
  wire g_59_55;
  wire p_59_56;
  wire g_59_56;
  wire p_59_57;
  wire g_59_57;
  wire p_59_58;
  wire g_59_58;
  wire p_60_60;
  wire g_60_60;
 assign p_60_60 = a[60] ^ b[60];
 assign g_60_60 = a[60] & b[60];
  wire p_60_0;
  wire g_60_0;
  wire p_60_1;
  wire g_60_1;
  wire p_60_2;
  wire g_60_2;
  wire p_60_3;
  wire g_60_3;
  wire p_60_4;
  wire g_60_4;
  wire p_60_5;
  wire g_60_5;
  wire p_60_6;
  wire g_60_6;
  wire p_60_7;
  wire g_60_7;
  wire p_60_8;
  wire g_60_8;
  wire p_60_9;
  wire g_60_9;
  wire p_60_10;
  wire g_60_10;
  wire p_60_11;
  wire g_60_11;
  wire p_60_12;
  wire g_60_12;
  wire p_60_13;
  wire g_60_13;
  wire p_60_14;
  wire g_60_14;
  wire p_60_15;
  wire g_60_15;
  wire p_60_16;
  wire g_60_16;
  wire p_60_17;
  wire g_60_17;
  wire p_60_18;
  wire g_60_18;
  wire p_60_19;
  wire g_60_19;
  wire p_60_20;
  wire g_60_20;
  wire p_60_21;
  wire g_60_21;
  wire p_60_22;
  wire g_60_22;
  wire p_60_23;
  wire g_60_23;
  wire p_60_24;
  wire g_60_24;
  wire p_60_25;
  wire g_60_25;
  wire p_60_26;
  wire g_60_26;
  wire p_60_27;
  wire g_60_27;
  wire p_60_28;
  wire g_60_28;
  wire p_60_29;
  wire g_60_29;
  wire p_60_30;
  wire g_60_30;
  wire p_60_31;
  wire g_60_31;
  wire p_60_32;
  wire g_60_32;
  wire p_60_33;
  wire g_60_33;
  wire p_60_34;
  wire g_60_34;
  wire p_60_35;
  wire g_60_35;
  wire p_60_36;
  wire g_60_36;
  wire p_60_37;
  wire g_60_37;
  wire p_60_38;
  wire g_60_38;
  wire p_60_39;
  wire g_60_39;
  wire p_60_40;
  wire g_60_40;
  wire p_60_41;
  wire g_60_41;
  wire p_60_42;
  wire g_60_42;
  wire p_60_43;
  wire g_60_43;
  wire p_60_44;
  wire g_60_44;
  wire p_60_45;
  wire g_60_45;
  wire p_60_46;
  wire g_60_46;
  wire p_60_47;
  wire g_60_47;
  wire p_60_48;
  wire g_60_48;
  wire p_60_49;
  wire g_60_49;
  wire p_60_50;
  wire g_60_50;
  wire p_60_51;
  wire g_60_51;
  wire p_60_52;
  wire g_60_52;
  wire p_60_53;
  wire g_60_53;
  wire p_60_54;
  wire g_60_54;
  wire p_60_55;
  wire g_60_55;
  wire p_60_56;
  wire g_60_56;
  wire p_60_57;
  wire g_60_57;
  wire p_60_58;
  wire g_60_58;
  wire p_60_59;
  wire g_60_59;
  wire p_61_61;
  wire g_61_61;
 assign p_61_61 = a[61] ^ b[61];
 assign g_61_61 = a[61] & b[61];
  wire p_61_0;
  wire g_61_0;
  wire p_61_1;
  wire g_61_1;
  wire p_61_2;
  wire g_61_2;
  wire p_61_3;
  wire g_61_3;
  wire p_61_4;
  wire g_61_4;
  wire p_61_5;
  wire g_61_5;
  wire p_61_6;
  wire g_61_6;
  wire p_61_7;
  wire g_61_7;
  wire p_61_8;
  wire g_61_8;
  wire p_61_9;
  wire g_61_9;
  wire p_61_10;
  wire g_61_10;
  wire p_61_11;
  wire g_61_11;
  wire p_61_12;
  wire g_61_12;
  wire p_61_13;
  wire g_61_13;
  wire p_61_14;
  wire g_61_14;
  wire p_61_15;
  wire g_61_15;
  wire p_61_16;
  wire g_61_16;
  wire p_61_17;
  wire g_61_17;
  wire p_61_18;
  wire g_61_18;
  wire p_61_19;
  wire g_61_19;
  wire p_61_20;
  wire g_61_20;
  wire p_61_21;
  wire g_61_21;
  wire p_61_22;
  wire g_61_22;
  wire p_61_23;
  wire g_61_23;
  wire p_61_24;
  wire g_61_24;
  wire p_61_25;
  wire g_61_25;
  wire p_61_26;
  wire g_61_26;
  wire p_61_27;
  wire g_61_27;
  wire p_61_28;
  wire g_61_28;
  wire p_61_29;
  wire g_61_29;
  wire p_61_30;
  wire g_61_30;
  wire p_61_31;
  wire g_61_31;
  wire p_61_32;
  wire g_61_32;
  wire p_61_33;
  wire g_61_33;
  wire p_61_34;
  wire g_61_34;
  wire p_61_35;
  wire g_61_35;
  wire p_61_36;
  wire g_61_36;
  wire p_61_37;
  wire g_61_37;
  wire p_61_38;
  wire g_61_38;
  wire p_61_39;
  wire g_61_39;
  wire p_61_40;
  wire g_61_40;
  wire p_61_41;
  wire g_61_41;
  wire p_61_42;
  wire g_61_42;
  wire p_61_43;
  wire g_61_43;
  wire p_61_44;
  wire g_61_44;
  wire p_61_45;
  wire g_61_45;
  wire p_61_46;
  wire g_61_46;
  wire p_61_47;
  wire g_61_47;
  wire p_61_48;
  wire g_61_48;
  wire p_61_49;
  wire g_61_49;
  wire p_61_50;
  wire g_61_50;
  wire p_61_51;
  wire g_61_51;
  wire p_61_52;
  wire g_61_52;
  wire p_61_53;
  wire g_61_53;
  wire p_61_54;
  wire g_61_54;
  wire p_61_55;
  wire g_61_55;
  wire p_61_56;
  wire g_61_56;
  wire p_61_57;
  wire g_61_57;
  wire p_61_58;
  wire g_61_58;
  wire p_61_59;
  wire g_61_59;
  wire p_61_60;
  wire g_61_60;
  wire p_62_62;
  wire g_62_62;
 assign p_62_62 = a[62] ^ b[62];
 assign g_62_62 = a[62] & b[62];
  wire p_62_0;
  wire g_62_0;
  wire p_62_1;
  wire g_62_1;
  wire p_62_2;
  wire g_62_2;
  wire p_62_3;
  wire g_62_3;
  wire p_62_4;
  wire g_62_4;
  wire p_62_5;
  wire g_62_5;
  wire p_62_6;
  wire g_62_6;
  wire p_62_7;
  wire g_62_7;
  wire p_62_8;
  wire g_62_8;
  wire p_62_9;
  wire g_62_9;
  wire p_62_10;
  wire g_62_10;
  wire p_62_11;
  wire g_62_11;
  wire p_62_12;
  wire g_62_12;
  wire p_62_13;
  wire g_62_13;
  wire p_62_14;
  wire g_62_14;
  wire p_62_15;
  wire g_62_15;
  wire p_62_16;
  wire g_62_16;
  wire p_62_17;
  wire g_62_17;
  wire p_62_18;
  wire g_62_18;
  wire p_62_19;
  wire g_62_19;
  wire p_62_20;
  wire g_62_20;
  wire p_62_21;
  wire g_62_21;
  wire p_62_22;
  wire g_62_22;
  wire p_62_23;
  wire g_62_23;
  wire p_62_24;
  wire g_62_24;
  wire p_62_25;
  wire g_62_25;
  wire p_62_26;
  wire g_62_26;
  wire p_62_27;
  wire g_62_27;
  wire p_62_28;
  wire g_62_28;
  wire p_62_29;
  wire g_62_29;
  wire p_62_30;
  wire g_62_30;
  wire p_62_31;
  wire g_62_31;
  wire p_62_32;
  wire g_62_32;
  wire p_62_33;
  wire g_62_33;
  wire p_62_34;
  wire g_62_34;
  wire p_62_35;
  wire g_62_35;
  wire p_62_36;
  wire g_62_36;
  wire p_62_37;
  wire g_62_37;
  wire p_62_38;
  wire g_62_38;
  wire p_62_39;
  wire g_62_39;
  wire p_62_40;
  wire g_62_40;
  wire p_62_41;
  wire g_62_41;
  wire p_62_42;
  wire g_62_42;
  wire p_62_43;
  wire g_62_43;
  wire p_62_44;
  wire g_62_44;
  wire p_62_45;
  wire g_62_45;
  wire p_62_46;
  wire g_62_46;
  wire p_62_47;
  wire g_62_47;
  wire p_62_48;
  wire g_62_48;
  wire p_62_49;
  wire g_62_49;
  wire p_62_50;
  wire g_62_50;
  wire p_62_51;
  wire g_62_51;
  wire p_62_52;
  wire g_62_52;
  wire p_62_53;
  wire g_62_53;
  wire p_62_54;
  wire g_62_54;
  wire p_62_55;
  wire g_62_55;
  wire p_62_56;
  wire g_62_56;
  wire p_62_57;
  wire g_62_57;
  wire p_62_58;
  wire g_62_58;
  wire p_62_59;
  wire g_62_59;
  wire p_62_60;
  wire g_62_60;
  wire p_62_61;
  wire g_62_61;
 assign sum[0] = p_0_0;
 assign p_1_0 = p_1_1 & p_0_0;
 assign g_1_0 = g_1_1 | (p_1_1 & g_0_0);
 assign sum[1] = p_1_1^ g_0_0;
 assign p_2_0 = p_2_1 & p_0_0;
 assign g_2_0 = g_2_1 | (p_2_1 & g_0_0);
 assign p_2_1 = p_2_2 & p_1_1;
 assign g_2_1 = g_2_2 | (p_2_2 & g_1_1);
 assign sum[2] = p_2_2^ g_1_0;
 assign p_3_0 = p_3_2 & p_1_0;
 assign g_3_0 = g_3_2 | (p_3_2 & g_1_0);
 assign p_3_1 = p_3_2 & p_1_1;
 assign g_3_1 = g_3_2 | (p_3_2 & g_1_1);
 assign p_3_2 = p_3_3 & p_2_2;
 assign g_3_2 = g_3_3 | (p_3_3 & g_2_2);
 assign sum[3] = p_3_3^ g_2_0;
 assign p_4_0 = p_4_1 & p_0_0;
 assign g_4_0 = g_4_1 | (p_4_1 & g_0_0);
 assign p_4_1 = p_4_3 & p_2_1;
 assign g_4_1 = g_4_3 | (p_4_3 & g_2_1);
 assign p_4_2 = p_4_3 & p_2_2;
 assign g_4_2 = g_4_3 | (p_4_3 & g_2_2);
 assign p_4_3 = p_4_4 & p_3_3;
 assign g_4_3 = g_4_4 | (p_4_4 & g_3_3);
 assign sum[4] = p_4_4^ g_3_0;
 assign p_5_0 = p_5_2 & p_1_0;
 assign g_5_0 = g_5_2 | (p_5_2 & g_1_0);
 assign p_5_1 = p_5_2 & p_1_1;
 assign g_5_1 = g_5_2 | (p_5_2 & g_1_1);
 assign p_5_2 = p_5_4 & p_3_2;
 assign g_5_2 = g_5_4 | (p_5_4 & g_3_2);
 assign p_5_3 = p_5_4 & p_3_3;
 assign g_5_3 = g_5_4 | (p_5_4 & g_3_3);
 assign p_5_4 = p_5_5 & p_4_4;
 assign g_5_4 = g_5_5 | (p_5_5 & g_4_4);
 assign sum[5] = p_5_5^ g_4_0;
 assign p_6_0 = p_6_3 & p_2_0;
 assign g_6_0 = g_6_3 | (p_6_3 & g_2_0);
 assign p_6_1 = p_6_3 & p_2_1;
 assign g_6_1 = g_6_3 | (p_6_3 & g_2_1);
 assign p_6_2 = p_6_3 & p_2_2;
 assign g_6_2 = g_6_3 | (p_6_3 & g_2_2);
 assign p_6_3 = p_6_5 & p_4_3;
 assign g_6_3 = g_6_5 | (p_6_5 & g_4_3);
 assign p_6_4 = p_6_5 & p_4_4;
 assign g_6_4 = g_6_5 | (p_6_5 & g_4_4);
 assign p_6_5 = p_6_6 & p_5_5;
 assign g_6_5 = g_6_6 | (p_6_6 & g_5_5);
 assign sum[6] = p_6_6^ g_5_0;
 assign p_7_0 = p_7_4 & p_3_0;
 assign g_7_0 = g_7_4 | (p_7_4 & g_3_0);
 assign p_7_1 = p_7_4 & p_3_1;
 assign g_7_1 = g_7_4 | (p_7_4 & g_3_1);
 assign p_7_2 = p_7_4 & p_3_2;
 assign g_7_2 = g_7_4 | (p_7_4 & g_3_2);
 assign p_7_3 = p_7_4 & p_3_3;
 assign g_7_3 = g_7_4 | (p_7_4 & g_3_3);
 assign p_7_4 = p_7_6 & p_5_4;
 assign g_7_4 = g_7_6 | (p_7_6 & g_5_4);
 assign p_7_5 = p_7_6 & p_5_5;
 assign g_7_5 = g_7_6 | (p_7_6 & g_5_5);
 assign p_7_6 = p_7_7 & p_6_6;
 assign g_7_6 = g_7_7 | (p_7_7 & g_6_6);
 assign sum[7] = p_7_7^ g_6_0;
 assign p_8_0 = p_8_1 & p_0_0;
 assign g_8_0 = g_8_1 | (p_8_1 & g_0_0);
 assign p_8_1 = p_8_5 & p_4_1;
 assign g_8_1 = g_8_5 | (p_8_5 & g_4_1);
 assign p_8_2 = p_8_5 & p_4_2;
 assign g_8_2 = g_8_5 | (p_8_5 & g_4_2);
 assign p_8_3 = p_8_5 & p_4_3;
 assign g_8_3 = g_8_5 | (p_8_5 & g_4_3);
 assign p_8_4 = p_8_5 & p_4_4;
 assign g_8_4 = g_8_5 | (p_8_5 & g_4_4);
 assign p_8_5 = p_8_7 & p_6_5;
 assign g_8_5 = g_8_7 | (p_8_7 & g_6_5);
 assign p_8_6 = p_8_7 & p_6_6;
 assign g_8_6 = g_8_7 | (p_8_7 & g_6_6);
 assign p_8_7 = p_8_8 & p_7_7;
 assign g_8_7 = g_8_8 | (p_8_8 & g_7_7);
 assign sum[8] = p_8_8^ g_7_0;
 assign p_9_0 = p_9_2 & p_1_0;
 assign g_9_0 = g_9_2 | (p_9_2 & g_1_0);
 assign p_9_1 = p_9_2 & p_1_1;
 assign g_9_1 = g_9_2 | (p_9_2 & g_1_1);
 assign p_9_2 = p_9_6 & p_5_2;
 assign g_9_2 = g_9_6 | (p_9_6 & g_5_2);
 assign p_9_3 = p_9_6 & p_5_3;
 assign g_9_3 = g_9_6 | (p_9_6 & g_5_3);
 assign p_9_4 = p_9_6 & p_5_4;
 assign g_9_4 = g_9_6 | (p_9_6 & g_5_4);
 assign p_9_5 = p_9_6 & p_5_5;
 assign g_9_5 = g_9_6 | (p_9_6 & g_5_5);
 assign p_9_6 = p_9_8 & p_7_6;
 assign g_9_6 = g_9_8 | (p_9_8 & g_7_6);
 assign p_9_7 = p_9_8 & p_7_7;
 assign g_9_7 = g_9_8 | (p_9_8 & g_7_7);
 assign p_9_8 = p_9_9 & p_8_8;
 assign g_9_8 = g_9_9 | (p_9_9 & g_8_8);
 assign sum[9] = p_9_9^ g_8_0;
 assign p_10_0 = p_10_3 & p_2_0;
 assign g_10_0 = g_10_3 | (p_10_3 & g_2_0);
 assign p_10_1 = p_10_3 & p_2_1;
 assign g_10_1 = g_10_3 | (p_10_3 & g_2_1);
 assign p_10_2 = p_10_3 & p_2_2;
 assign g_10_2 = g_10_3 | (p_10_3 & g_2_2);
 assign p_10_3 = p_10_7 & p_6_3;
 assign g_10_3 = g_10_7 | (p_10_7 & g_6_3);
 assign p_10_4 = p_10_7 & p_6_4;
 assign g_10_4 = g_10_7 | (p_10_7 & g_6_4);
 assign p_10_5 = p_10_7 & p_6_5;
 assign g_10_5 = g_10_7 | (p_10_7 & g_6_5);
 assign p_10_6 = p_10_7 & p_6_6;
 assign g_10_6 = g_10_7 | (p_10_7 & g_6_6);
 assign p_10_7 = p_10_9 & p_8_7;
 assign g_10_7 = g_10_9 | (p_10_9 & g_8_7);
 assign p_10_8 = p_10_9 & p_8_8;
 assign g_10_8 = g_10_9 | (p_10_9 & g_8_8);
 assign p_10_9 = p_10_10 & p_9_9;
 assign g_10_9 = g_10_10 | (p_10_10 & g_9_9);
 assign sum[10] = p_10_10^ g_9_0;
 assign p_11_0 = p_11_4 & p_3_0;
 assign g_11_0 = g_11_4 | (p_11_4 & g_3_0);
 assign p_11_1 = p_11_4 & p_3_1;
 assign g_11_1 = g_11_4 | (p_11_4 & g_3_1);
 assign p_11_2 = p_11_4 & p_3_2;
 assign g_11_2 = g_11_4 | (p_11_4 & g_3_2);
 assign p_11_3 = p_11_4 & p_3_3;
 assign g_11_3 = g_11_4 | (p_11_4 & g_3_3);
 assign p_11_4 = p_11_8 & p_7_4;
 assign g_11_4 = g_11_8 | (p_11_8 & g_7_4);
 assign p_11_5 = p_11_8 & p_7_5;
 assign g_11_5 = g_11_8 | (p_11_8 & g_7_5);
 assign p_11_6 = p_11_8 & p_7_6;
 assign g_11_6 = g_11_8 | (p_11_8 & g_7_6);
 assign p_11_7 = p_11_8 & p_7_7;
 assign g_11_7 = g_11_8 | (p_11_8 & g_7_7);
 assign p_11_8 = p_11_10 & p_9_8;
 assign g_11_8 = g_11_10 | (p_11_10 & g_9_8);
 assign p_11_9 = p_11_10 & p_9_9;
 assign g_11_9 = g_11_10 | (p_11_10 & g_9_9);
 assign p_11_10 = p_11_11 & p_10_10;
 assign g_11_10 = g_11_11 | (p_11_11 & g_10_10);
 assign sum[11] = p_11_11^ g_10_0;
 assign p_12_0 = p_12_5 & p_4_0;
 assign g_12_0 = g_12_5 | (p_12_5 & g_4_0);
 assign p_12_1 = p_12_5 & p_4_1;
 assign g_12_1 = g_12_5 | (p_12_5 & g_4_1);
 assign p_12_2 = p_12_5 & p_4_2;
 assign g_12_2 = g_12_5 | (p_12_5 & g_4_2);
 assign p_12_3 = p_12_5 & p_4_3;
 assign g_12_3 = g_12_5 | (p_12_5 & g_4_3);
 assign p_12_4 = p_12_5 & p_4_4;
 assign g_12_4 = g_12_5 | (p_12_5 & g_4_4);
 assign p_12_5 = p_12_9 & p_8_5;
 assign g_12_5 = g_12_9 | (p_12_9 & g_8_5);
 assign p_12_6 = p_12_9 & p_8_6;
 assign g_12_6 = g_12_9 | (p_12_9 & g_8_6);
 assign p_12_7 = p_12_9 & p_8_7;
 assign g_12_7 = g_12_9 | (p_12_9 & g_8_7);
 assign p_12_8 = p_12_9 & p_8_8;
 assign g_12_8 = g_12_9 | (p_12_9 & g_8_8);
 assign p_12_9 = p_12_11 & p_10_9;
 assign g_12_9 = g_12_11 | (p_12_11 & g_10_9);
 assign p_12_10 = p_12_11 & p_10_10;
 assign g_12_10 = g_12_11 | (p_12_11 & g_10_10);
 assign p_12_11 = p_12_12 & p_11_11;
 assign g_12_11 = g_12_12 | (p_12_12 & g_11_11);
 assign sum[12] = p_12_12^ g_11_0;
 assign p_13_0 = p_13_6 & p_5_0;
 assign g_13_0 = g_13_6 | (p_13_6 & g_5_0);
 assign p_13_1 = p_13_6 & p_5_1;
 assign g_13_1 = g_13_6 | (p_13_6 & g_5_1);
 assign p_13_2 = p_13_6 & p_5_2;
 assign g_13_2 = g_13_6 | (p_13_6 & g_5_2);
 assign p_13_3 = p_13_6 & p_5_3;
 assign g_13_3 = g_13_6 | (p_13_6 & g_5_3);
 assign p_13_4 = p_13_6 & p_5_4;
 assign g_13_4 = g_13_6 | (p_13_6 & g_5_4);
 assign p_13_5 = p_13_6 & p_5_5;
 assign g_13_5 = g_13_6 | (p_13_6 & g_5_5);
 assign p_13_6 = p_13_10 & p_9_6;
 assign g_13_6 = g_13_10 | (p_13_10 & g_9_6);
 assign p_13_7 = p_13_10 & p_9_7;
 assign g_13_7 = g_13_10 | (p_13_10 & g_9_7);
 assign p_13_8 = p_13_10 & p_9_8;
 assign g_13_8 = g_13_10 | (p_13_10 & g_9_8);
 assign p_13_9 = p_13_10 & p_9_9;
 assign g_13_9 = g_13_10 | (p_13_10 & g_9_9);
 assign p_13_10 = p_13_12 & p_11_10;
 assign g_13_10 = g_13_12 | (p_13_12 & g_11_10);
 assign p_13_11 = p_13_12 & p_11_11;
 assign g_13_11 = g_13_12 | (p_13_12 & g_11_11);
 assign p_13_12 = p_13_13 & p_12_12;
 assign g_13_12 = g_13_13 | (p_13_13 & g_12_12);
 assign sum[13] = p_13_13^ g_12_0;
 assign p_14_0 = p_14_7 & p_6_0;
 assign g_14_0 = g_14_7 | (p_14_7 & g_6_0);
 assign p_14_1 = p_14_7 & p_6_1;
 assign g_14_1 = g_14_7 | (p_14_7 & g_6_1);
 assign p_14_2 = p_14_7 & p_6_2;
 assign g_14_2 = g_14_7 | (p_14_7 & g_6_2);
 assign p_14_3 = p_14_7 & p_6_3;
 assign g_14_3 = g_14_7 | (p_14_7 & g_6_3);
 assign p_14_4 = p_14_7 & p_6_4;
 assign g_14_4 = g_14_7 | (p_14_7 & g_6_4);
 assign p_14_5 = p_14_7 & p_6_5;
 assign g_14_5 = g_14_7 | (p_14_7 & g_6_5);
 assign p_14_6 = p_14_7 & p_6_6;
 assign g_14_6 = g_14_7 | (p_14_7 & g_6_6);
 assign p_14_7 = p_14_11 & p_10_7;
 assign g_14_7 = g_14_11 | (p_14_11 & g_10_7);
 assign p_14_8 = p_14_11 & p_10_8;
 assign g_14_8 = g_14_11 | (p_14_11 & g_10_8);
 assign p_14_9 = p_14_11 & p_10_9;
 assign g_14_9 = g_14_11 | (p_14_11 & g_10_9);
 assign p_14_10 = p_14_11 & p_10_10;
 assign g_14_10 = g_14_11 | (p_14_11 & g_10_10);
 assign p_14_11 = p_14_13 & p_12_11;
 assign g_14_11 = g_14_13 | (p_14_13 & g_12_11);
 assign p_14_12 = p_14_13 & p_12_12;
 assign g_14_12 = g_14_13 | (p_14_13 & g_12_12);
 assign p_14_13 = p_14_14 & p_13_13;
 assign g_14_13 = g_14_14 | (p_14_14 & g_13_13);
 assign sum[14] = p_14_14^ g_13_0;
 assign p_15_0 = p_15_8 & p_7_0;
 assign g_15_0 = g_15_8 | (p_15_8 & g_7_0);
 assign p_15_1 = p_15_8 & p_7_1;
 assign g_15_1 = g_15_8 | (p_15_8 & g_7_1);
 assign p_15_2 = p_15_8 & p_7_2;
 assign g_15_2 = g_15_8 | (p_15_8 & g_7_2);
 assign p_15_3 = p_15_8 & p_7_3;
 assign g_15_3 = g_15_8 | (p_15_8 & g_7_3);
 assign p_15_4 = p_15_8 & p_7_4;
 assign g_15_4 = g_15_8 | (p_15_8 & g_7_4);
 assign p_15_5 = p_15_8 & p_7_5;
 assign g_15_5 = g_15_8 | (p_15_8 & g_7_5);
 assign p_15_6 = p_15_8 & p_7_6;
 assign g_15_6 = g_15_8 | (p_15_8 & g_7_6);
 assign p_15_7 = p_15_8 & p_7_7;
 assign g_15_7 = g_15_8 | (p_15_8 & g_7_7);
 assign p_15_8 = p_15_12 & p_11_8;
 assign g_15_8 = g_15_12 | (p_15_12 & g_11_8);
 assign p_15_9 = p_15_12 & p_11_9;
 assign g_15_9 = g_15_12 | (p_15_12 & g_11_9);
 assign p_15_10 = p_15_12 & p_11_10;
 assign g_15_10 = g_15_12 | (p_15_12 & g_11_10);
 assign p_15_11 = p_15_12 & p_11_11;
 assign g_15_11 = g_15_12 | (p_15_12 & g_11_11);
 assign p_15_12 = p_15_14 & p_13_12;
 assign g_15_12 = g_15_14 | (p_15_14 & g_13_12);
 assign p_15_13 = p_15_14 & p_13_13;
 assign g_15_13 = g_15_14 | (p_15_14 & g_13_13);
 assign p_15_14 = p_15_15 & p_14_14;
 assign g_15_14 = g_15_15 | (p_15_15 & g_14_14);
 assign sum[15] = p_15_15^ g_14_0;
 assign p_16_0 = p_16_1 & p_0_0;
 assign g_16_0 = g_16_1 | (p_16_1 & g_0_0);
 assign p_16_1 = p_16_9 & p_8_1;
 assign g_16_1 = g_16_9 | (p_16_9 & g_8_1);
 assign p_16_2 = p_16_9 & p_8_2;
 assign g_16_2 = g_16_9 | (p_16_9 & g_8_2);
 assign p_16_3 = p_16_9 & p_8_3;
 assign g_16_3 = g_16_9 | (p_16_9 & g_8_3);
 assign p_16_4 = p_16_9 & p_8_4;
 assign g_16_4 = g_16_9 | (p_16_9 & g_8_4);
 assign p_16_5 = p_16_9 & p_8_5;
 assign g_16_5 = g_16_9 | (p_16_9 & g_8_5);
 assign p_16_6 = p_16_9 & p_8_6;
 assign g_16_6 = g_16_9 | (p_16_9 & g_8_6);
 assign p_16_7 = p_16_9 & p_8_7;
 assign g_16_7 = g_16_9 | (p_16_9 & g_8_7);
 assign p_16_8 = p_16_9 & p_8_8;
 assign g_16_8 = g_16_9 | (p_16_9 & g_8_8);
 assign p_16_9 = p_16_13 & p_12_9;
 assign g_16_9 = g_16_13 | (p_16_13 & g_12_9);
 assign p_16_10 = p_16_13 & p_12_10;
 assign g_16_10 = g_16_13 | (p_16_13 & g_12_10);
 assign p_16_11 = p_16_13 & p_12_11;
 assign g_16_11 = g_16_13 | (p_16_13 & g_12_11);
 assign p_16_12 = p_16_13 & p_12_12;
 assign g_16_12 = g_16_13 | (p_16_13 & g_12_12);
 assign p_16_13 = p_16_15 & p_14_13;
 assign g_16_13 = g_16_15 | (p_16_15 & g_14_13);
 assign p_16_14 = p_16_15 & p_14_14;
 assign g_16_14 = g_16_15 | (p_16_15 & g_14_14);
 assign p_16_15 = p_16_16 & p_15_15;
 assign g_16_15 = g_16_16 | (p_16_16 & g_15_15);
 assign sum[16] = p_16_16^ g_15_0;
 assign p_17_0 = p_17_2 & p_1_0;
 assign g_17_0 = g_17_2 | (p_17_2 & g_1_0);
 assign p_17_1 = p_17_2 & p_1_1;
 assign g_17_1 = g_17_2 | (p_17_2 & g_1_1);
 assign p_17_2 = p_17_10 & p_9_2;
 assign g_17_2 = g_17_10 | (p_17_10 & g_9_2);
 assign p_17_3 = p_17_10 & p_9_3;
 assign g_17_3 = g_17_10 | (p_17_10 & g_9_3);
 assign p_17_4 = p_17_10 & p_9_4;
 assign g_17_4 = g_17_10 | (p_17_10 & g_9_4);
 assign p_17_5 = p_17_10 & p_9_5;
 assign g_17_5 = g_17_10 | (p_17_10 & g_9_5);
 assign p_17_6 = p_17_10 & p_9_6;
 assign g_17_6 = g_17_10 | (p_17_10 & g_9_6);
 assign p_17_7 = p_17_10 & p_9_7;
 assign g_17_7 = g_17_10 | (p_17_10 & g_9_7);
 assign p_17_8 = p_17_10 & p_9_8;
 assign g_17_8 = g_17_10 | (p_17_10 & g_9_8);
 assign p_17_9 = p_17_10 & p_9_9;
 assign g_17_9 = g_17_10 | (p_17_10 & g_9_9);
 assign p_17_10 = p_17_14 & p_13_10;
 assign g_17_10 = g_17_14 | (p_17_14 & g_13_10);
 assign p_17_11 = p_17_14 & p_13_11;
 assign g_17_11 = g_17_14 | (p_17_14 & g_13_11);
 assign p_17_12 = p_17_14 & p_13_12;
 assign g_17_12 = g_17_14 | (p_17_14 & g_13_12);
 assign p_17_13 = p_17_14 & p_13_13;
 assign g_17_13 = g_17_14 | (p_17_14 & g_13_13);
 assign p_17_14 = p_17_16 & p_15_14;
 assign g_17_14 = g_17_16 | (p_17_16 & g_15_14);
 assign p_17_15 = p_17_16 & p_15_15;
 assign g_17_15 = g_17_16 | (p_17_16 & g_15_15);
 assign p_17_16 = p_17_17 & p_16_16;
 assign g_17_16 = g_17_17 | (p_17_17 & g_16_16);
 assign sum[17] = p_17_17^ g_16_0;
 assign p_18_0 = p_18_3 & p_2_0;
 assign g_18_0 = g_18_3 | (p_18_3 & g_2_0);
 assign p_18_1 = p_18_3 & p_2_1;
 assign g_18_1 = g_18_3 | (p_18_3 & g_2_1);
 assign p_18_2 = p_18_3 & p_2_2;
 assign g_18_2 = g_18_3 | (p_18_3 & g_2_2);
 assign p_18_3 = p_18_11 & p_10_3;
 assign g_18_3 = g_18_11 | (p_18_11 & g_10_3);
 assign p_18_4 = p_18_11 & p_10_4;
 assign g_18_4 = g_18_11 | (p_18_11 & g_10_4);
 assign p_18_5 = p_18_11 & p_10_5;
 assign g_18_5 = g_18_11 | (p_18_11 & g_10_5);
 assign p_18_6 = p_18_11 & p_10_6;
 assign g_18_6 = g_18_11 | (p_18_11 & g_10_6);
 assign p_18_7 = p_18_11 & p_10_7;
 assign g_18_7 = g_18_11 | (p_18_11 & g_10_7);
 assign p_18_8 = p_18_11 & p_10_8;
 assign g_18_8 = g_18_11 | (p_18_11 & g_10_8);
 assign p_18_9 = p_18_11 & p_10_9;
 assign g_18_9 = g_18_11 | (p_18_11 & g_10_9);
 assign p_18_10 = p_18_11 & p_10_10;
 assign g_18_10 = g_18_11 | (p_18_11 & g_10_10);
 assign p_18_11 = p_18_15 & p_14_11;
 assign g_18_11 = g_18_15 | (p_18_15 & g_14_11);
 assign p_18_12 = p_18_15 & p_14_12;
 assign g_18_12 = g_18_15 | (p_18_15 & g_14_12);
 assign p_18_13 = p_18_15 & p_14_13;
 assign g_18_13 = g_18_15 | (p_18_15 & g_14_13);
 assign p_18_14 = p_18_15 & p_14_14;
 assign g_18_14 = g_18_15 | (p_18_15 & g_14_14);
 assign p_18_15 = p_18_17 & p_16_15;
 assign g_18_15 = g_18_17 | (p_18_17 & g_16_15);
 assign p_18_16 = p_18_17 & p_16_16;
 assign g_18_16 = g_18_17 | (p_18_17 & g_16_16);
 assign p_18_17 = p_18_18 & p_17_17;
 assign g_18_17 = g_18_18 | (p_18_18 & g_17_17);
 assign sum[18] = p_18_18^ g_17_0;
 assign p_19_0 = p_19_4 & p_3_0;
 assign g_19_0 = g_19_4 | (p_19_4 & g_3_0);
 assign p_19_1 = p_19_4 & p_3_1;
 assign g_19_1 = g_19_4 | (p_19_4 & g_3_1);
 assign p_19_2 = p_19_4 & p_3_2;
 assign g_19_2 = g_19_4 | (p_19_4 & g_3_2);
 assign p_19_3 = p_19_4 & p_3_3;
 assign g_19_3 = g_19_4 | (p_19_4 & g_3_3);
 assign p_19_4 = p_19_12 & p_11_4;
 assign g_19_4 = g_19_12 | (p_19_12 & g_11_4);
 assign p_19_5 = p_19_12 & p_11_5;
 assign g_19_5 = g_19_12 | (p_19_12 & g_11_5);
 assign p_19_6 = p_19_12 & p_11_6;
 assign g_19_6 = g_19_12 | (p_19_12 & g_11_6);
 assign p_19_7 = p_19_12 & p_11_7;
 assign g_19_7 = g_19_12 | (p_19_12 & g_11_7);
 assign p_19_8 = p_19_12 & p_11_8;
 assign g_19_8 = g_19_12 | (p_19_12 & g_11_8);
 assign p_19_9 = p_19_12 & p_11_9;
 assign g_19_9 = g_19_12 | (p_19_12 & g_11_9);
 assign p_19_10 = p_19_12 & p_11_10;
 assign g_19_10 = g_19_12 | (p_19_12 & g_11_10);
 assign p_19_11 = p_19_12 & p_11_11;
 assign g_19_11 = g_19_12 | (p_19_12 & g_11_11);
 assign p_19_12 = p_19_16 & p_15_12;
 assign g_19_12 = g_19_16 | (p_19_16 & g_15_12);
 assign p_19_13 = p_19_16 & p_15_13;
 assign g_19_13 = g_19_16 | (p_19_16 & g_15_13);
 assign p_19_14 = p_19_16 & p_15_14;
 assign g_19_14 = g_19_16 | (p_19_16 & g_15_14);
 assign p_19_15 = p_19_16 & p_15_15;
 assign g_19_15 = g_19_16 | (p_19_16 & g_15_15);
 assign p_19_16 = p_19_18 & p_17_16;
 assign g_19_16 = g_19_18 | (p_19_18 & g_17_16);
 assign p_19_17 = p_19_18 & p_17_17;
 assign g_19_17 = g_19_18 | (p_19_18 & g_17_17);
 assign p_19_18 = p_19_19 & p_18_18;
 assign g_19_18 = g_19_19 | (p_19_19 & g_18_18);
 assign sum[19] = p_19_19^ g_18_0;
 assign p_20_0 = p_20_5 & p_4_0;
 assign g_20_0 = g_20_5 | (p_20_5 & g_4_0);
 assign p_20_1 = p_20_5 & p_4_1;
 assign g_20_1 = g_20_5 | (p_20_5 & g_4_1);
 assign p_20_2 = p_20_5 & p_4_2;
 assign g_20_2 = g_20_5 | (p_20_5 & g_4_2);
 assign p_20_3 = p_20_5 & p_4_3;
 assign g_20_3 = g_20_5 | (p_20_5 & g_4_3);
 assign p_20_4 = p_20_5 & p_4_4;
 assign g_20_4 = g_20_5 | (p_20_5 & g_4_4);
 assign p_20_5 = p_20_13 & p_12_5;
 assign g_20_5 = g_20_13 | (p_20_13 & g_12_5);
 assign p_20_6 = p_20_13 & p_12_6;
 assign g_20_6 = g_20_13 | (p_20_13 & g_12_6);
 assign p_20_7 = p_20_13 & p_12_7;
 assign g_20_7 = g_20_13 | (p_20_13 & g_12_7);
 assign p_20_8 = p_20_13 & p_12_8;
 assign g_20_8 = g_20_13 | (p_20_13 & g_12_8);
 assign p_20_9 = p_20_13 & p_12_9;
 assign g_20_9 = g_20_13 | (p_20_13 & g_12_9);
 assign p_20_10 = p_20_13 & p_12_10;
 assign g_20_10 = g_20_13 | (p_20_13 & g_12_10);
 assign p_20_11 = p_20_13 & p_12_11;
 assign g_20_11 = g_20_13 | (p_20_13 & g_12_11);
 assign p_20_12 = p_20_13 & p_12_12;
 assign g_20_12 = g_20_13 | (p_20_13 & g_12_12);
 assign p_20_13 = p_20_17 & p_16_13;
 assign g_20_13 = g_20_17 | (p_20_17 & g_16_13);
 assign p_20_14 = p_20_17 & p_16_14;
 assign g_20_14 = g_20_17 | (p_20_17 & g_16_14);
 assign p_20_15 = p_20_17 & p_16_15;
 assign g_20_15 = g_20_17 | (p_20_17 & g_16_15);
 assign p_20_16 = p_20_17 & p_16_16;
 assign g_20_16 = g_20_17 | (p_20_17 & g_16_16);
 assign p_20_17 = p_20_19 & p_18_17;
 assign g_20_17 = g_20_19 | (p_20_19 & g_18_17);
 assign p_20_18 = p_20_19 & p_18_18;
 assign g_20_18 = g_20_19 | (p_20_19 & g_18_18);
 assign p_20_19 = p_20_20 & p_19_19;
 assign g_20_19 = g_20_20 | (p_20_20 & g_19_19);
 assign sum[20] = p_20_20^ g_19_0;
 assign p_21_0 = p_21_6 & p_5_0;
 assign g_21_0 = g_21_6 | (p_21_6 & g_5_0);
 assign p_21_1 = p_21_6 & p_5_1;
 assign g_21_1 = g_21_6 | (p_21_6 & g_5_1);
 assign p_21_2 = p_21_6 & p_5_2;
 assign g_21_2 = g_21_6 | (p_21_6 & g_5_2);
 assign p_21_3 = p_21_6 & p_5_3;
 assign g_21_3 = g_21_6 | (p_21_6 & g_5_3);
 assign p_21_4 = p_21_6 & p_5_4;
 assign g_21_4 = g_21_6 | (p_21_6 & g_5_4);
 assign p_21_5 = p_21_6 & p_5_5;
 assign g_21_5 = g_21_6 | (p_21_6 & g_5_5);
 assign p_21_6 = p_21_14 & p_13_6;
 assign g_21_6 = g_21_14 | (p_21_14 & g_13_6);
 assign p_21_7 = p_21_14 & p_13_7;
 assign g_21_7 = g_21_14 | (p_21_14 & g_13_7);
 assign p_21_8 = p_21_14 & p_13_8;
 assign g_21_8 = g_21_14 | (p_21_14 & g_13_8);
 assign p_21_9 = p_21_14 & p_13_9;
 assign g_21_9 = g_21_14 | (p_21_14 & g_13_9);
 assign p_21_10 = p_21_14 & p_13_10;
 assign g_21_10 = g_21_14 | (p_21_14 & g_13_10);
 assign p_21_11 = p_21_14 & p_13_11;
 assign g_21_11 = g_21_14 | (p_21_14 & g_13_11);
 assign p_21_12 = p_21_14 & p_13_12;
 assign g_21_12 = g_21_14 | (p_21_14 & g_13_12);
 assign p_21_13 = p_21_14 & p_13_13;
 assign g_21_13 = g_21_14 | (p_21_14 & g_13_13);
 assign p_21_14 = p_21_18 & p_17_14;
 assign g_21_14 = g_21_18 | (p_21_18 & g_17_14);
 assign p_21_15 = p_21_18 & p_17_15;
 assign g_21_15 = g_21_18 | (p_21_18 & g_17_15);
 assign p_21_16 = p_21_18 & p_17_16;
 assign g_21_16 = g_21_18 | (p_21_18 & g_17_16);
 assign p_21_17 = p_21_18 & p_17_17;
 assign g_21_17 = g_21_18 | (p_21_18 & g_17_17);
 assign p_21_18 = p_21_20 & p_19_18;
 assign g_21_18 = g_21_20 | (p_21_20 & g_19_18);
 assign p_21_19 = p_21_20 & p_19_19;
 assign g_21_19 = g_21_20 | (p_21_20 & g_19_19);
 assign p_21_20 = p_21_21 & p_20_20;
 assign g_21_20 = g_21_21 | (p_21_21 & g_20_20);
 assign sum[21] = p_21_21^ g_20_0;
 assign p_22_0 = p_22_7 & p_6_0;
 assign g_22_0 = g_22_7 | (p_22_7 & g_6_0);
 assign p_22_1 = p_22_7 & p_6_1;
 assign g_22_1 = g_22_7 | (p_22_7 & g_6_1);
 assign p_22_2 = p_22_7 & p_6_2;
 assign g_22_2 = g_22_7 | (p_22_7 & g_6_2);
 assign p_22_3 = p_22_7 & p_6_3;
 assign g_22_3 = g_22_7 | (p_22_7 & g_6_3);
 assign p_22_4 = p_22_7 & p_6_4;
 assign g_22_4 = g_22_7 | (p_22_7 & g_6_4);
 assign p_22_5 = p_22_7 & p_6_5;
 assign g_22_5 = g_22_7 | (p_22_7 & g_6_5);
 assign p_22_6 = p_22_7 & p_6_6;
 assign g_22_6 = g_22_7 | (p_22_7 & g_6_6);
 assign p_22_7 = p_22_15 & p_14_7;
 assign g_22_7 = g_22_15 | (p_22_15 & g_14_7);
 assign p_22_8 = p_22_15 & p_14_8;
 assign g_22_8 = g_22_15 | (p_22_15 & g_14_8);
 assign p_22_9 = p_22_15 & p_14_9;
 assign g_22_9 = g_22_15 | (p_22_15 & g_14_9);
 assign p_22_10 = p_22_15 & p_14_10;
 assign g_22_10 = g_22_15 | (p_22_15 & g_14_10);
 assign p_22_11 = p_22_15 & p_14_11;
 assign g_22_11 = g_22_15 | (p_22_15 & g_14_11);
 assign p_22_12 = p_22_15 & p_14_12;
 assign g_22_12 = g_22_15 | (p_22_15 & g_14_12);
 assign p_22_13 = p_22_15 & p_14_13;
 assign g_22_13 = g_22_15 | (p_22_15 & g_14_13);
 assign p_22_14 = p_22_15 & p_14_14;
 assign g_22_14 = g_22_15 | (p_22_15 & g_14_14);
 assign p_22_15 = p_22_19 & p_18_15;
 assign g_22_15 = g_22_19 | (p_22_19 & g_18_15);
 assign p_22_16 = p_22_19 & p_18_16;
 assign g_22_16 = g_22_19 | (p_22_19 & g_18_16);
 assign p_22_17 = p_22_19 & p_18_17;
 assign g_22_17 = g_22_19 | (p_22_19 & g_18_17);
 assign p_22_18 = p_22_19 & p_18_18;
 assign g_22_18 = g_22_19 | (p_22_19 & g_18_18);
 assign p_22_19 = p_22_21 & p_20_19;
 assign g_22_19 = g_22_21 | (p_22_21 & g_20_19);
 assign p_22_20 = p_22_21 & p_20_20;
 assign g_22_20 = g_22_21 | (p_22_21 & g_20_20);
 assign p_22_21 = p_22_22 & p_21_21;
 assign g_22_21 = g_22_22 | (p_22_22 & g_21_21);
 assign sum[22] = p_22_22^ g_21_0;
 assign p_23_0 = p_23_8 & p_7_0;
 assign g_23_0 = g_23_8 | (p_23_8 & g_7_0);
 assign p_23_1 = p_23_8 & p_7_1;
 assign g_23_1 = g_23_8 | (p_23_8 & g_7_1);
 assign p_23_2 = p_23_8 & p_7_2;
 assign g_23_2 = g_23_8 | (p_23_8 & g_7_2);
 assign p_23_3 = p_23_8 & p_7_3;
 assign g_23_3 = g_23_8 | (p_23_8 & g_7_3);
 assign p_23_4 = p_23_8 & p_7_4;
 assign g_23_4 = g_23_8 | (p_23_8 & g_7_4);
 assign p_23_5 = p_23_8 & p_7_5;
 assign g_23_5 = g_23_8 | (p_23_8 & g_7_5);
 assign p_23_6 = p_23_8 & p_7_6;
 assign g_23_6 = g_23_8 | (p_23_8 & g_7_6);
 assign p_23_7 = p_23_8 & p_7_7;
 assign g_23_7 = g_23_8 | (p_23_8 & g_7_7);
 assign p_23_8 = p_23_16 & p_15_8;
 assign g_23_8 = g_23_16 | (p_23_16 & g_15_8);
 assign p_23_9 = p_23_16 & p_15_9;
 assign g_23_9 = g_23_16 | (p_23_16 & g_15_9);
 assign p_23_10 = p_23_16 & p_15_10;
 assign g_23_10 = g_23_16 | (p_23_16 & g_15_10);
 assign p_23_11 = p_23_16 & p_15_11;
 assign g_23_11 = g_23_16 | (p_23_16 & g_15_11);
 assign p_23_12 = p_23_16 & p_15_12;
 assign g_23_12 = g_23_16 | (p_23_16 & g_15_12);
 assign p_23_13 = p_23_16 & p_15_13;
 assign g_23_13 = g_23_16 | (p_23_16 & g_15_13);
 assign p_23_14 = p_23_16 & p_15_14;
 assign g_23_14 = g_23_16 | (p_23_16 & g_15_14);
 assign p_23_15 = p_23_16 & p_15_15;
 assign g_23_15 = g_23_16 | (p_23_16 & g_15_15);
 assign p_23_16 = p_23_20 & p_19_16;
 assign g_23_16 = g_23_20 | (p_23_20 & g_19_16);
 assign p_23_17 = p_23_20 & p_19_17;
 assign g_23_17 = g_23_20 | (p_23_20 & g_19_17);
 assign p_23_18 = p_23_20 & p_19_18;
 assign g_23_18 = g_23_20 | (p_23_20 & g_19_18);
 assign p_23_19 = p_23_20 & p_19_19;
 assign g_23_19 = g_23_20 | (p_23_20 & g_19_19);
 assign p_23_20 = p_23_22 & p_21_20;
 assign g_23_20 = g_23_22 | (p_23_22 & g_21_20);
 assign p_23_21 = p_23_22 & p_21_21;
 assign g_23_21 = g_23_22 | (p_23_22 & g_21_21);
 assign p_23_22 = p_23_23 & p_22_22;
 assign g_23_22 = g_23_23 | (p_23_23 & g_22_22);
 assign sum[23] = p_23_23^ g_22_0;
 assign p_24_0 = p_24_9 & p_8_0;
 assign g_24_0 = g_24_9 | (p_24_9 & g_8_0);
 assign p_24_1 = p_24_9 & p_8_1;
 assign g_24_1 = g_24_9 | (p_24_9 & g_8_1);
 assign p_24_2 = p_24_9 & p_8_2;
 assign g_24_2 = g_24_9 | (p_24_9 & g_8_2);
 assign p_24_3 = p_24_9 & p_8_3;
 assign g_24_3 = g_24_9 | (p_24_9 & g_8_3);
 assign p_24_4 = p_24_9 & p_8_4;
 assign g_24_4 = g_24_9 | (p_24_9 & g_8_4);
 assign p_24_5 = p_24_9 & p_8_5;
 assign g_24_5 = g_24_9 | (p_24_9 & g_8_5);
 assign p_24_6 = p_24_9 & p_8_6;
 assign g_24_6 = g_24_9 | (p_24_9 & g_8_6);
 assign p_24_7 = p_24_9 & p_8_7;
 assign g_24_7 = g_24_9 | (p_24_9 & g_8_7);
 assign p_24_8 = p_24_9 & p_8_8;
 assign g_24_8 = g_24_9 | (p_24_9 & g_8_8);
 assign p_24_9 = p_24_17 & p_16_9;
 assign g_24_9 = g_24_17 | (p_24_17 & g_16_9);
 assign p_24_10 = p_24_17 & p_16_10;
 assign g_24_10 = g_24_17 | (p_24_17 & g_16_10);
 assign p_24_11 = p_24_17 & p_16_11;
 assign g_24_11 = g_24_17 | (p_24_17 & g_16_11);
 assign p_24_12 = p_24_17 & p_16_12;
 assign g_24_12 = g_24_17 | (p_24_17 & g_16_12);
 assign p_24_13 = p_24_17 & p_16_13;
 assign g_24_13 = g_24_17 | (p_24_17 & g_16_13);
 assign p_24_14 = p_24_17 & p_16_14;
 assign g_24_14 = g_24_17 | (p_24_17 & g_16_14);
 assign p_24_15 = p_24_17 & p_16_15;
 assign g_24_15 = g_24_17 | (p_24_17 & g_16_15);
 assign p_24_16 = p_24_17 & p_16_16;
 assign g_24_16 = g_24_17 | (p_24_17 & g_16_16);
 assign p_24_17 = p_24_21 & p_20_17;
 assign g_24_17 = g_24_21 | (p_24_21 & g_20_17);
 assign p_24_18 = p_24_21 & p_20_18;
 assign g_24_18 = g_24_21 | (p_24_21 & g_20_18);
 assign p_24_19 = p_24_21 & p_20_19;
 assign g_24_19 = g_24_21 | (p_24_21 & g_20_19);
 assign p_24_20 = p_24_21 & p_20_20;
 assign g_24_20 = g_24_21 | (p_24_21 & g_20_20);
 assign p_24_21 = p_24_23 & p_22_21;
 assign g_24_21 = g_24_23 | (p_24_23 & g_22_21);
 assign p_24_22 = p_24_23 & p_22_22;
 assign g_24_22 = g_24_23 | (p_24_23 & g_22_22);
 assign p_24_23 = p_24_24 & p_23_23;
 assign g_24_23 = g_24_24 | (p_24_24 & g_23_23);
 assign sum[24] = p_24_24^ g_23_0;
 assign p_25_0 = p_25_10 & p_9_0;
 assign g_25_0 = g_25_10 | (p_25_10 & g_9_0);
 assign p_25_1 = p_25_10 & p_9_1;
 assign g_25_1 = g_25_10 | (p_25_10 & g_9_1);
 assign p_25_2 = p_25_10 & p_9_2;
 assign g_25_2 = g_25_10 | (p_25_10 & g_9_2);
 assign p_25_3 = p_25_10 & p_9_3;
 assign g_25_3 = g_25_10 | (p_25_10 & g_9_3);
 assign p_25_4 = p_25_10 & p_9_4;
 assign g_25_4 = g_25_10 | (p_25_10 & g_9_4);
 assign p_25_5 = p_25_10 & p_9_5;
 assign g_25_5 = g_25_10 | (p_25_10 & g_9_5);
 assign p_25_6 = p_25_10 & p_9_6;
 assign g_25_6 = g_25_10 | (p_25_10 & g_9_6);
 assign p_25_7 = p_25_10 & p_9_7;
 assign g_25_7 = g_25_10 | (p_25_10 & g_9_7);
 assign p_25_8 = p_25_10 & p_9_8;
 assign g_25_8 = g_25_10 | (p_25_10 & g_9_8);
 assign p_25_9 = p_25_10 & p_9_9;
 assign g_25_9 = g_25_10 | (p_25_10 & g_9_9);
 assign p_25_10 = p_25_18 & p_17_10;
 assign g_25_10 = g_25_18 | (p_25_18 & g_17_10);
 assign p_25_11 = p_25_18 & p_17_11;
 assign g_25_11 = g_25_18 | (p_25_18 & g_17_11);
 assign p_25_12 = p_25_18 & p_17_12;
 assign g_25_12 = g_25_18 | (p_25_18 & g_17_12);
 assign p_25_13 = p_25_18 & p_17_13;
 assign g_25_13 = g_25_18 | (p_25_18 & g_17_13);
 assign p_25_14 = p_25_18 & p_17_14;
 assign g_25_14 = g_25_18 | (p_25_18 & g_17_14);
 assign p_25_15 = p_25_18 & p_17_15;
 assign g_25_15 = g_25_18 | (p_25_18 & g_17_15);
 assign p_25_16 = p_25_18 & p_17_16;
 assign g_25_16 = g_25_18 | (p_25_18 & g_17_16);
 assign p_25_17 = p_25_18 & p_17_17;
 assign g_25_17 = g_25_18 | (p_25_18 & g_17_17);
 assign p_25_18 = p_25_22 & p_21_18;
 assign g_25_18 = g_25_22 | (p_25_22 & g_21_18);
 assign p_25_19 = p_25_22 & p_21_19;
 assign g_25_19 = g_25_22 | (p_25_22 & g_21_19);
 assign p_25_20 = p_25_22 & p_21_20;
 assign g_25_20 = g_25_22 | (p_25_22 & g_21_20);
 assign p_25_21 = p_25_22 & p_21_21;
 assign g_25_21 = g_25_22 | (p_25_22 & g_21_21);
 assign p_25_22 = p_25_24 & p_23_22;
 assign g_25_22 = g_25_24 | (p_25_24 & g_23_22);
 assign p_25_23 = p_25_24 & p_23_23;
 assign g_25_23 = g_25_24 | (p_25_24 & g_23_23);
 assign p_25_24 = p_25_25 & p_24_24;
 assign g_25_24 = g_25_25 | (p_25_25 & g_24_24);
 assign sum[25] = p_25_25^ g_24_0;
 assign p_26_0 = p_26_11 & p_10_0;
 assign g_26_0 = g_26_11 | (p_26_11 & g_10_0);
 assign p_26_1 = p_26_11 & p_10_1;
 assign g_26_1 = g_26_11 | (p_26_11 & g_10_1);
 assign p_26_2 = p_26_11 & p_10_2;
 assign g_26_2 = g_26_11 | (p_26_11 & g_10_2);
 assign p_26_3 = p_26_11 & p_10_3;
 assign g_26_3 = g_26_11 | (p_26_11 & g_10_3);
 assign p_26_4 = p_26_11 & p_10_4;
 assign g_26_4 = g_26_11 | (p_26_11 & g_10_4);
 assign p_26_5 = p_26_11 & p_10_5;
 assign g_26_5 = g_26_11 | (p_26_11 & g_10_5);
 assign p_26_6 = p_26_11 & p_10_6;
 assign g_26_6 = g_26_11 | (p_26_11 & g_10_6);
 assign p_26_7 = p_26_11 & p_10_7;
 assign g_26_7 = g_26_11 | (p_26_11 & g_10_7);
 assign p_26_8 = p_26_11 & p_10_8;
 assign g_26_8 = g_26_11 | (p_26_11 & g_10_8);
 assign p_26_9 = p_26_11 & p_10_9;
 assign g_26_9 = g_26_11 | (p_26_11 & g_10_9);
 assign p_26_10 = p_26_11 & p_10_10;
 assign g_26_10 = g_26_11 | (p_26_11 & g_10_10);
 assign p_26_11 = p_26_19 & p_18_11;
 assign g_26_11 = g_26_19 | (p_26_19 & g_18_11);
 assign p_26_12 = p_26_19 & p_18_12;
 assign g_26_12 = g_26_19 | (p_26_19 & g_18_12);
 assign p_26_13 = p_26_19 & p_18_13;
 assign g_26_13 = g_26_19 | (p_26_19 & g_18_13);
 assign p_26_14 = p_26_19 & p_18_14;
 assign g_26_14 = g_26_19 | (p_26_19 & g_18_14);
 assign p_26_15 = p_26_19 & p_18_15;
 assign g_26_15 = g_26_19 | (p_26_19 & g_18_15);
 assign p_26_16 = p_26_19 & p_18_16;
 assign g_26_16 = g_26_19 | (p_26_19 & g_18_16);
 assign p_26_17 = p_26_19 & p_18_17;
 assign g_26_17 = g_26_19 | (p_26_19 & g_18_17);
 assign p_26_18 = p_26_19 & p_18_18;
 assign g_26_18 = g_26_19 | (p_26_19 & g_18_18);
 assign p_26_19 = p_26_23 & p_22_19;
 assign g_26_19 = g_26_23 | (p_26_23 & g_22_19);
 assign p_26_20 = p_26_23 & p_22_20;
 assign g_26_20 = g_26_23 | (p_26_23 & g_22_20);
 assign p_26_21 = p_26_23 & p_22_21;
 assign g_26_21 = g_26_23 | (p_26_23 & g_22_21);
 assign p_26_22 = p_26_23 & p_22_22;
 assign g_26_22 = g_26_23 | (p_26_23 & g_22_22);
 assign p_26_23 = p_26_25 & p_24_23;
 assign g_26_23 = g_26_25 | (p_26_25 & g_24_23);
 assign p_26_24 = p_26_25 & p_24_24;
 assign g_26_24 = g_26_25 | (p_26_25 & g_24_24);
 assign p_26_25 = p_26_26 & p_25_25;
 assign g_26_25 = g_26_26 | (p_26_26 & g_25_25);
 assign sum[26] = p_26_26^ g_25_0;
 assign p_27_0 = p_27_12 & p_11_0;
 assign g_27_0 = g_27_12 | (p_27_12 & g_11_0);
 assign p_27_1 = p_27_12 & p_11_1;
 assign g_27_1 = g_27_12 | (p_27_12 & g_11_1);
 assign p_27_2 = p_27_12 & p_11_2;
 assign g_27_2 = g_27_12 | (p_27_12 & g_11_2);
 assign p_27_3 = p_27_12 & p_11_3;
 assign g_27_3 = g_27_12 | (p_27_12 & g_11_3);
 assign p_27_4 = p_27_12 & p_11_4;
 assign g_27_4 = g_27_12 | (p_27_12 & g_11_4);
 assign p_27_5 = p_27_12 & p_11_5;
 assign g_27_5 = g_27_12 | (p_27_12 & g_11_5);
 assign p_27_6 = p_27_12 & p_11_6;
 assign g_27_6 = g_27_12 | (p_27_12 & g_11_6);
 assign p_27_7 = p_27_12 & p_11_7;
 assign g_27_7 = g_27_12 | (p_27_12 & g_11_7);
 assign p_27_8 = p_27_12 & p_11_8;
 assign g_27_8 = g_27_12 | (p_27_12 & g_11_8);
 assign p_27_9 = p_27_12 & p_11_9;
 assign g_27_9 = g_27_12 | (p_27_12 & g_11_9);
 assign p_27_10 = p_27_12 & p_11_10;
 assign g_27_10 = g_27_12 | (p_27_12 & g_11_10);
 assign p_27_11 = p_27_12 & p_11_11;
 assign g_27_11 = g_27_12 | (p_27_12 & g_11_11);
 assign p_27_12 = p_27_20 & p_19_12;
 assign g_27_12 = g_27_20 | (p_27_20 & g_19_12);
 assign p_27_13 = p_27_20 & p_19_13;
 assign g_27_13 = g_27_20 | (p_27_20 & g_19_13);
 assign p_27_14 = p_27_20 & p_19_14;
 assign g_27_14 = g_27_20 | (p_27_20 & g_19_14);
 assign p_27_15 = p_27_20 & p_19_15;
 assign g_27_15 = g_27_20 | (p_27_20 & g_19_15);
 assign p_27_16 = p_27_20 & p_19_16;
 assign g_27_16 = g_27_20 | (p_27_20 & g_19_16);
 assign p_27_17 = p_27_20 & p_19_17;
 assign g_27_17 = g_27_20 | (p_27_20 & g_19_17);
 assign p_27_18 = p_27_20 & p_19_18;
 assign g_27_18 = g_27_20 | (p_27_20 & g_19_18);
 assign p_27_19 = p_27_20 & p_19_19;
 assign g_27_19 = g_27_20 | (p_27_20 & g_19_19);
 assign p_27_20 = p_27_24 & p_23_20;
 assign g_27_20 = g_27_24 | (p_27_24 & g_23_20);
 assign p_27_21 = p_27_24 & p_23_21;
 assign g_27_21 = g_27_24 | (p_27_24 & g_23_21);
 assign p_27_22 = p_27_24 & p_23_22;
 assign g_27_22 = g_27_24 | (p_27_24 & g_23_22);
 assign p_27_23 = p_27_24 & p_23_23;
 assign g_27_23 = g_27_24 | (p_27_24 & g_23_23);
 assign p_27_24 = p_27_26 & p_25_24;
 assign g_27_24 = g_27_26 | (p_27_26 & g_25_24);
 assign p_27_25 = p_27_26 & p_25_25;
 assign g_27_25 = g_27_26 | (p_27_26 & g_25_25);
 assign p_27_26 = p_27_27 & p_26_26;
 assign g_27_26 = g_27_27 | (p_27_27 & g_26_26);
 assign sum[27] = p_27_27^ g_26_0;
 assign p_28_0 = p_28_13 & p_12_0;
 assign g_28_0 = g_28_13 | (p_28_13 & g_12_0);
 assign p_28_1 = p_28_13 & p_12_1;
 assign g_28_1 = g_28_13 | (p_28_13 & g_12_1);
 assign p_28_2 = p_28_13 & p_12_2;
 assign g_28_2 = g_28_13 | (p_28_13 & g_12_2);
 assign p_28_3 = p_28_13 & p_12_3;
 assign g_28_3 = g_28_13 | (p_28_13 & g_12_3);
 assign p_28_4 = p_28_13 & p_12_4;
 assign g_28_4 = g_28_13 | (p_28_13 & g_12_4);
 assign p_28_5 = p_28_13 & p_12_5;
 assign g_28_5 = g_28_13 | (p_28_13 & g_12_5);
 assign p_28_6 = p_28_13 & p_12_6;
 assign g_28_6 = g_28_13 | (p_28_13 & g_12_6);
 assign p_28_7 = p_28_13 & p_12_7;
 assign g_28_7 = g_28_13 | (p_28_13 & g_12_7);
 assign p_28_8 = p_28_13 & p_12_8;
 assign g_28_8 = g_28_13 | (p_28_13 & g_12_8);
 assign p_28_9 = p_28_13 & p_12_9;
 assign g_28_9 = g_28_13 | (p_28_13 & g_12_9);
 assign p_28_10 = p_28_13 & p_12_10;
 assign g_28_10 = g_28_13 | (p_28_13 & g_12_10);
 assign p_28_11 = p_28_13 & p_12_11;
 assign g_28_11 = g_28_13 | (p_28_13 & g_12_11);
 assign p_28_12 = p_28_13 & p_12_12;
 assign g_28_12 = g_28_13 | (p_28_13 & g_12_12);
 assign p_28_13 = p_28_21 & p_20_13;
 assign g_28_13 = g_28_21 | (p_28_21 & g_20_13);
 assign p_28_14 = p_28_21 & p_20_14;
 assign g_28_14 = g_28_21 | (p_28_21 & g_20_14);
 assign p_28_15 = p_28_21 & p_20_15;
 assign g_28_15 = g_28_21 | (p_28_21 & g_20_15);
 assign p_28_16 = p_28_21 & p_20_16;
 assign g_28_16 = g_28_21 | (p_28_21 & g_20_16);
 assign p_28_17 = p_28_21 & p_20_17;
 assign g_28_17 = g_28_21 | (p_28_21 & g_20_17);
 assign p_28_18 = p_28_21 & p_20_18;
 assign g_28_18 = g_28_21 | (p_28_21 & g_20_18);
 assign p_28_19 = p_28_21 & p_20_19;
 assign g_28_19 = g_28_21 | (p_28_21 & g_20_19);
 assign p_28_20 = p_28_21 & p_20_20;
 assign g_28_20 = g_28_21 | (p_28_21 & g_20_20);
 assign p_28_21 = p_28_25 & p_24_21;
 assign g_28_21 = g_28_25 | (p_28_25 & g_24_21);
 assign p_28_22 = p_28_25 & p_24_22;
 assign g_28_22 = g_28_25 | (p_28_25 & g_24_22);
 assign p_28_23 = p_28_25 & p_24_23;
 assign g_28_23 = g_28_25 | (p_28_25 & g_24_23);
 assign p_28_24 = p_28_25 & p_24_24;
 assign g_28_24 = g_28_25 | (p_28_25 & g_24_24);
 assign p_28_25 = p_28_27 & p_26_25;
 assign g_28_25 = g_28_27 | (p_28_27 & g_26_25);
 assign p_28_26 = p_28_27 & p_26_26;
 assign g_28_26 = g_28_27 | (p_28_27 & g_26_26);
 assign p_28_27 = p_28_28 & p_27_27;
 assign g_28_27 = g_28_28 | (p_28_28 & g_27_27);
 assign sum[28] = p_28_28^ g_27_0;
 assign p_29_0 = p_29_14 & p_13_0;
 assign g_29_0 = g_29_14 | (p_29_14 & g_13_0);
 assign p_29_1 = p_29_14 & p_13_1;
 assign g_29_1 = g_29_14 | (p_29_14 & g_13_1);
 assign p_29_2 = p_29_14 & p_13_2;
 assign g_29_2 = g_29_14 | (p_29_14 & g_13_2);
 assign p_29_3 = p_29_14 & p_13_3;
 assign g_29_3 = g_29_14 | (p_29_14 & g_13_3);
 assign p_29_4 = p_29_14 & p_13_4;
 assign g_29_4 = g_29_14 | (p_29_14 & g_13_4);
 assign p_29_5 = p_29_14 & p_13_5;
 assign g_29_5 = g_29_14 | (p_29_14 & g_13_5);
 assign p_29_6 = p_29_14 & p_13_6;
 assign g_29_6 = g_29_14 | (p_29_14 & g_13_6);
 assign p_29_7 = p_29_14 & p_13_7;
 assign g_29_7 = g_29_14 | (p_29_14 & g_13_7);
 assign p_29_8 = p_29_14 & p_13_8;
 assign g_29_8 = g_29_14 | (p_29_14 & g_13_8);
 assign p_29_9 = p_29_14 & p_13_9;
 assign g_29_9 = g_29_14 | (p_29_14 & g_13_9);
 assign p_29_10 = p_29_14 & p_13_10;
 assign g_29_10 = g_29_14 | (p_29_14 & g_13_10);
 assign p_29_11 = p_29_14 & p_13_11;
 assign g_29_11 = g_29_14 | (p_29_14 & g_13_11);
 assign p_29_12 = p_29_14 & p_13_12;
 assign g_29_12 = g_29_14 | (p_29_14 & g_13_12);
 assign p_29_13 = p_29_14 & p_13_13;
 assign g_29_13 = g_29_14 | (p_29_14 & g_13_13);
 assign p_29_14 = p_29_22 & p_21_14;
 assign g_29_14 = g_29_22 | (p_29_22 & g_21_14);
 assign p_29_15 = p_29_22 & p_21_15;
 assign g_29_15 = g_29_22 | (p_29_22 & g_21_15);
 assign p_29_16 = p_29_22 & p_21_16;
 assign g_29_16 = g_29_22 | (p_29_22 & g_21_16);
 assign p_29_17 = p_29_22 & p_21_17;
 assign g_29_17 = g_29_22 | (p_29_22 & g_21_17);
 assign p_29_18 = p_29_22 & p_21_18;
 assign g_29_18 = g_29_22 | (p_29_22 & g_21_18);
 assign p_29_19 = p_29_22 & p_21_19;
 assign g_29_19 = g_29_22 | (p_29_22 & g_21_19);
 assign p_29_20 = p_29_22 & p_21_20;
 assign g_29_20 = g_29_22 | (p_29_22 & g_21_20);
 assign p_29_21 = p_29_22 & p_21_21;
 assign g_29_21 = g_29_22 | (p_29_22 & g_21_21);
 assign p_29_22 = p_29_26 & p_25_22;
 assign g_29_22 = g_29_26 | (p_29_26 & g_25_22);
 assign p_29_23 = p_29_26 & p_25_23;
 assign g_29_23 = g_29_26 | (p_29_26 & g_25_23);
 assign p_29_24 = p_29_26 & p_25_24;
 assign g_29_24 = g_29_26 | (p_29_26 & g_25_24);
 assign p_29_25 = p_29_26 & p_25_25;
 assign g_29_25 = g_29_26 | (p_29_26 & g_25_25);
 assign p_29_26 = p_29_28 & p_27_26;
 assign g_29_26 = g_29_28 | (p_29_28 & g_27_26);
 assign p_29_27 = p_29_28 & p_27_27;
 assign g_29_27 = g_29_28 | (p_29_28 & g_27_27);
 assign p_29_28 = p_29_29 & p_28_28;
 assign g_29_28 = g_29_29 | (p_29_29 & g_28_28);
 assign sum[29] = p_29_29^ g_28_0;
 assign p_30_0 = p_30_15 & p_14_0;
 assign g_30_0 = g_30_15 | (p_30_15 & g_14_0);
 assign p_30_1 = p_30_15 & p_14_1;
 assign g_30_1 = g_30_15 | (p_30_15 & g_14_1);
 assign p_30_2 = p_30_15 & p_14_2;
 assign g_30_2 = g_30_15 | (p_30_15 & g_14_2);
 assign p_30_3 = p_30_15 & p_14_3;
 assign g_30_3 = g_30_15 | (p_30_15 & g_14_3);
 assign p_30_4 = p_30_15 & p_14_4;
 assign g_30_4 = g_30_15 | (p_30_15 & g_14_4);
 assign p_30_5 = p_30_15 & p_14_5;
 assign g_30_5 = g_30_15 | (p_30_15 & g_14_5);
 assign p_30_6 = p_30_15 & p_14_6;
 assign g_30_6 = g_30_15 | (p_30_15 & g_14_6);
 assign p_30_7 = p_30_15 & p_14_7;
 assign g_30_7 = g_30_15 | (p_30_15 & g_14_7);
 assign p_30_8 = p_30_15 & p_14_8;
 assign g_30_8 = g_30_15 | (p_30_15 & g_14_8);
 assign p_30_9 = p_30_15 & p_14_9;
 assign g_30_9 = g_30_15 | (p_30_15 & g_14_9);
 assign p_30_10 = p_30_15 & p_14_10;
 assign g_30_10 = g_30_15 | (p_30_15 & g_14_10);
 assign p_30_11 = p_30_15 & p_14_11;
 assign g_30_11 = g_30_15 | (p_30_15 & g_14_11);
 assign p_30_12 = p_30_15 & p_14_12;
 assign g_30_12 = g_30_15 | (p_30_15 & g_14_12);
 assign p_30_13 = p_30_15 & p_14_13;
 assign g_30_13 = g_30_15 | (p_30_15 & g_14_13);
 assign p_30_14 = p_30_15 & p_14_14;
 assign g_30_14 = g_30_15 | (p_30_15 & g_14_14);
 assign p_30_15 = p_30_23 & p_22_15;
 assign g_30_15 = g_30_23 | (p_30_23 & g_22_15);
 assign p_30_16 = p_30_23 & p_22_16;
 assign g_30_16 = g_30_23 | (p_30_23 & g_22_16);
 assign p_30_17 = p_30_23 & p_22_17;
 assign g_30_17 = g_30_23 | (p_30_23 & g_22_17);
 assign p_30_18 = p_30_23 & p_22_18;
 assign g_30_18 = g_30_23 | (p_30_23 & g_22_18);
 assign p_30_19 = p_30_23 & p_22_19;
 assign g_30_19 = g_30_23 | (p_30_23 & g_22_19);
 assign p_30_20 = p_30_23 & p_22_20;
 assign g_30_20 = g_30_23 | (p_30_23 & g_22_20);
 assign p_30_21 = p_30_23 & p_22_21;
 assign g_30_21 = g_30_23 | (p_30_23 & g_22_21);
 assign p_30_22 = p_30_23 & p_22_22;
 assign g_30_22 = g_30_23 | (p_30_23 & g_22_22);
 assign p_30_23 = p_30_27 & p_26_23;
 assign g_30_23 = g_30_27 | (p_30_27 & g_26_23);
 assign p_30_24 = p_30_27 & p_26_24;
 assign g_30_24 = g_30_27 | (p_30_27 & g_26_24);
 assign p_30_25 = p_30_27 & p_26_25;
 assign g_30_25 = g_30_27 | (p_30_27 & g_26_25);
 assign p_30_26 = p_30_27 & p_26_26;
 assign g_30_26 = g_30_27 | (p_30_27 & g_26_26);
 assign p_30_27 = p_30_29 & p_28_27;
 assign g_30_27 = g_30_29 | (p_30_29 & g_28_27);
 assign p_30_28 = p_30_29 & p_28_28;
 assign g_30_28 = g_30_29 | (p_30_29 & g_28_28);
 assign p_30_29 = p_30_30 & p_29_29;
 assign g_30_29 = g_30_30 | (p_30_30 & g_29_29);
 assign sum[30] = p_30_30^ g_29_0;
 assign p_31_0 = p_31_16 & p_15_0;
 assign g_31_0 = g_31_16 | (p_31_16 & g_15_0);
 assign p_31_1 = p_31_16 & p_15_1;
 assign g_31_1 = g_31_16 | (p_31_16 & g_15_1);
 assign p_31_2 = p_31_16 & p_15_2;
 assign g_31_2 = g_31_16 | (p_31_16 & g_15_2);
 assign p_31_3 = p_31_16 & p_15_3;
 assign g_31_3 = g_31_16 | (p_31_16 & g_15_3);
 assign p_31_4 = p_31_16 & p_15_4;
 assign g_31_4 = g_31_16 | (p_31_16 & g_15_4);
 assign p_31_5 = p_31_16 & p_15_5;
 assign g_31_5 = g_31_16 | (p_31_16 & g_15_5);
 assign p_31_6 = p_31_16 & p_15_6;
 assign g_31_6 = g_31_16 | (p_31_16 & g_15_6);
 assign p_31_7 = p_31_16 & p_15_7;
 assign g_31_7 = g_31_16 | (p_31_16 & g_15_7);
 assign p_31_8 = p_31_16 & p_15_8;
 assign g_31_8 = g_31_16 | (p_31_16 & g_15_8);
 assign p_31_9 = p_31_16 & p_15_9;
 assign g_31_9 = g_31_16 | (p_31_16 & g_15_9);
 assign p_31_10 = p_31_16 & p_15_10;
 assign g_31_10 = g_31_16 | (p_31_16 & g_15_10);
 assign p_31_11 = p_31_16 & p_15_11;
 assign g_31_11 = g_31_16 | (p_31_16 & g_15_11);
 assign p_31_12 = p_31_16 & p_15_12;
 assign g_31_12 = g_31_16 | (p_31_16 & g_15_12);
 assign p_31_13 = p_31_16 & p_15_13;
 assign g_31_13 = g_31_16 | (p_31_16 & g_15_13);
 assign p_31_14 = p_31_16 & p_15_14;
 assign g_31_14 = g_31_16 | (p_31_16 & g_15_14);
 assign p_31_15 = p_31_16 & p_15_15;
 assign g_31_15 = g_31_16 | (p_31_16 & g_15_15);
 assign p_31_16 = p_31_24 & p_23_16;
 assign g_31_16 = g_31_24 | (p_31_24 & g_23_16);
 assign p_31_17 = p_31_24 & p_23_17;
 assign g_31_17 = g_31_24 | (p_31_24 & g_23_17);
 assign p_31_18 = p_31_24 & p_23_18;
 assign g_31_18 = g_31_24 | (p_31_24 & g_23_18);
 assign p_31_19 = p_31_24 & p_23_19;
 assign g_31_19 = g_31_24 | (p_31_24 & g_23_19);
 assign p_31_20 = p_31_24 & p_23_20;
 assign g_31_20 = g_31_24 | (p_31_24 & g_23_20);
 assign p_31_21 = p_31_24 & p_23_21;
 assign g_31_21 = g_31_24 | (p_31_24 & g_23_21);
 assign p_31_22 = p_31_24 & p_23_22;
 assign g_31_22 = g_31_24 | (p_31_24 & g_23_22);
 assign p_31_23 = p_31_24 & p_23_23;
 assign g_31_23 = g_31_24 | (p_31_24 & g_23_23);
 assign p_31_24 = p_31_28 & p_27_24;
 assign g_31_24 = g_31_28 | (p_31_28 & g_27_24);
 assign p_31_25 = p_31_28 & p_27_25;
 assign g_31_25 = g_31_28 | (p_31_28 & g_27_25);
 assign p_31_26 = p_31_28 & p_27_26;
 assign g_31_26 = g_31_28 | (p_31_28 & g_27_26);
 assign p_31_27 = p_31_28 & p_27_27;
 assign g_31_27 = g_31_28 | (p_31_28 & g_27_27);
 assign p_31_28 = p_31_30 & p_29_28;
 assign g_31_28 = g_31_30 | (p_31_30 & g_29_28);
 assign p_31_29 = p_31_30 & p_29_29;
 assign g_31_29 = g_31_30 | (p_31_30 & g_29_29);
 assign p_31_30 = p_31_31 & p_30_30;
 assign g_31_30 = g_31_31 | (p_31_31 & g_30_30);
 assign sum[31] = p_31_31^ g_30_0;
 assign p_32_0 = p_32_1 & p_0_0;
 assign g_32_0 = g_32_1 | (p_32_1 & g_0_0);
 assign p_32_1 = p_32_17 & p_16_1;
 assign g_32_1 = g_32_17 | (p_32_17 & g_16_1);
 assign p_32_2 = p_32_17 & p_16_2;
 assign g_32_2 = g_32_17 | (p_32_17 & g_16_2);
 assign p_32_3 = p_32_17 & p_16_3;
 assign g_32_3 = g_32_17 | (p_32_17 & g_16_3);
 assign p_32_4 = p_32_17 & p_16_4;
 assign g_32_4 = g_32_17 | (p_32_17 & g_16_4);
 assign p_32_5 = p_32_17 & p_16_5;
 assign g_32_5 = g_32_17 | (p_32_17 & g_16_5);
 assign p_32_6 = p_32_17 & p_16_6;
 assign g_32_6 = g_32_17 | (p_32_17 & g_16_6);
 assign p_32_7 = p_32_17 & p_16_7;
 assign g_32_7 = g_32_17 | (p_32_17 & g_16_7);
 assign p_32_8 = p_32_17 & p_16_8;
 assign g_32_8 = g_32_17 | (p_32_17 & g_16_8);
 assign p_32_9 = p_32_17 & p_16_9;
 assign g_32_9 = g_32_17 | (p_32_17 & g_16_9);
 assign p_32_10 = p_32_17 & p_16_10;
 assign g_32_10 = g_32_17 | (p_32_17 & g_16_10);
 assign p_32_11 = p_32_17 & p_16_11;
 assign g_32_11 = g_32_17 | (p_32_17 & g_16_11);
 assign p_32_12 = p_32_17 & p_16_12;
 assign g_32_12 = g_32_17 | (p_32_17 & g_16_12);
 assign p_32_13 = p_32_17 & p_16_13;
 assign g_32_13 = g_32_17 | (p_32_17 & g_16_13);
 assign p_32_14 = p_32_17 & p_16_14;
 assign g_32_14 = g_32_17 | (p_32_17 & g_16_14);
 assign p_32_15 = p_32_17 & p_16_15;
 assign g_32_15 = g_32_17 | (p_32_17 & g_16_15);
 assign p_32_16 = p_32_17 & p_16_16;
 assign g_32_16 = g_32_17 | (p_32_17 & g_16_16);
 assign p_32_17 = p_32_25 & p_24_17;
 assign g_32_17 = g_32_25 | (p_32_25 & g_24_17);
 assign p_32_18 = p_32_25 & p_24_18;
 assign g_32_18 = g_32_25 | (p_32_25 & g_24_18);
 assign p_32_19 = p_32_25 & p_24_19;
 assign g_32_19 = g_32_25 | (p_32_25 & g_24_19);
 assign p_32_20 = p_32_25 & p_24_20;
 assign g_32_20 = g_32_25 | (p_32_25 & g_24_20);
 assign p_32_21 = p_32_25 & p_24_21;
 assign g_32_21 = g_32_25 | (p_32_25 & g_24_21);
 assign p_32_22 = p_32_25 & p_24_22;
 assign g_32_22 = g_32_25 | (p_32_25 & g_24_22);
 assign p_32_23 = p_32_25 & p_24_23;
 assign g_32_23 = g_32_25 | (p_32_25 & g_24_23);
 assign p_32_24 = p_32_25 & p_24_24;
 assign g_32_24 = g_32_25 | (p_32_25 & g_24_24);
 assign p_32_25 = p_32_29 & p_28_25;
 assign g_32_25 = g_32_29 | (p_32_29 & g_28_25);
 assign p_32_26 = p_32_29 & p_28_26;
 assign g_32_26 = g_32_29 | (p_32_29 & g_28_26);
 assign p_32_27 = p_32_29 & p_28_27;
 assign g_32_27 = g_32_29 | (p_32_29 & g_28_27);
 assign p_32_28 = p_32_29 & p_28_28;
 assign g_32_28 = g_32_29 | (p_32_29 & g_28_28);
 assign p_32_29 = p_32_31 & p_30_29;
 assign g_32_29 = g_32_31 | (p_32_31 & g_30_29);
 assign p_32_30 = p_32_31 & p_30_30;
 assign g_32_30 = g_32_31 | (p_32_31 & g_30_30);
 assign p_32_31 = p_32_32 & p_31_31;
 assign g_32_31 = g_32_32 | (p_32_32 & g_31_31);
 assign sum[32] = p_32_32^ g_31_0;
 assign p_33_0 = p_33_2 & p_1_0;
 assign g_33_0 = g_33_2 | (p_33_2 & g_1_0);
 assign p_33_1 = p_33_2 & p_1_1;
 assign g_33_1 = g_33_2 | (p_33_2 & g_1_1);
 assign p_33_2 = p_33_18 & p_17_2;
 assign g_33_2 = g_33_18 | (p_33_18 & g_17_2);
 assign p_33_3 = p_33_18 & p_17_3;
 assign g_33_3 = g_33_18 | (p_33_18 & g_17_3);
 assign p_33_4 = p_33_18 & p_17_4;
 assign g_33_4 = g_33_18 | (p_33_18 & g_17_4);
 assign p_33_5 = p_33_18 & p_17_5;
 assign g_33_5 = g_33_18 | (p_33_18 & g_17_5);
 assign p_33_6 = p_33_18 & p_17_6;
 assign g_33_6 = g_33_18 | (p_33_18 & g_17_6);
 assign p_33_7 = p_33_18 & p_17_7;
 assign g_33_7 = g_33_18 | (p_33_18 & g_17_7);
 assign p_33_8 = p_33_18 & p_17_8;
 assign g_33_8 = g_33_18 | (p_33_18 & g_17_8);
 assign p_33_9 = p_33_18 & p_17_9;
 assign g_33_9 = g_33_18 | (p_33_18 & g_17_9);
 assign p_33_10 = p_33_18 & p_17_10;
 assign g_33_10 = g_33_18 | (p_33_18 & g_17_10);
 assign p_33_11 = p_33_18 & p_17_11;
 assign g_33_11 = g_33_18 | (p_33_18 & g_17_11);
 assign p_33_12 = p_33_18 & p_17_12;
 assign g_33_12 = g_33_18 | (p_33_18 & g_17_12);
 assign p_33_13 = p_33_18 & p_17_13;
 assign g_33_13 = g_33_18 | (p_33_18 & g_17_13);
 assign p_33_14 = p_33_18 & p_17_14;
 assign g_33_14 = g_33_18 | (p_33_18 & g_17_14);
 assign p_33_15 = p_33_18 & p_17_15;
 assign g_33_15 = g_33_18 | (p_33_18 & g_17_15);
 assign p_33_16 = p_33_18 & p_17_16;
 assign g_33_16 = g_33_18 | (p_33_18 & g_17_16);
 assign p_33_17 = p_33_18 & p_17_17;
 assign g_33_17 = g_33_18 | (p_33_18 & g_17_17);
 assign p_33_18 = p_33_26 & p_25_18;
 assign g_33_18 = g_33_26 | (p_33_26 & g_25_18);
 assign p_33_19 = p_33_26 & p_25_19;
 assign g_33_19 = g_33_26 | (p_33_26 & g_25_19);
 assign p_33_20 = p_33_26 & p_25_20;
 assign g_33_20 = g_33_26 | (p_33_26 & g_25_20);
 assign p_33_21 = p_33_26 & p_25_21;
 assign g_33_21 = g_33_26 | (p_33_26 & g_25_21);
 assign p_33_22 = p_33_26 & p_25_22;
 assign g_33_22 = g_33_26 | (p_33_26 & g_25_22);
 assign p_33_23 = p_33_26 & p_25_23;
 assign g_33_23 = g_33_26 | (p_33_26 & g_25_23);
 assign p_33_24 = p_33_26 & p_25_24;
 assign g_33_24 = g_33_26 | (p_33_26 & g_25_24);
 assign p_33_25 = p_33_26 & p_25_25;
 assign g_33_25 = g_33_26 | (p_33_26 & g_25_25);
 assign p_33_26 = p_33_30 & p_29_26;
 assign g_33_26 = g_33_30 | (p_33_30 & g_29_26);
 assign p_33_27 = p_33_30 & p_29_27;
 assign g_33_27 = g_33_30 | (p_33_30 & g_29_27);
 assign p_33_28 = p_33_30 & p_29_28;
 assign g_33_28 = g_33_30 | (p_33_30 & g_29_28);
 assign p_33_29 = p_33_30 & p_29_29;
 assign g_33_29 = g_33_30 | (p_33_30 & g_29_29);
 assign p_33_30 = p_33_32 & p_31_30;
 assign g_33_30 = g_33_32 | (p_33_32 & g_31_30);
 assign p_33_31 = p_33_32 & p_31_31;
 assign g_33_31 = g_33_32 | (p_33_32 & g_31_31);
 assign p_33_32 = p_33_33 & p_32_32;
 assign g_33_32 = g_33_33 | (p_33_33 & g_32_32);
 assign sum[33] = p_33_33^ g_32_0;
 assign p_34_0 = p_34_3 & p_2_0;
 assign g_34_0 = g_34_3 | (p_34_3 & g_2_0);
 assign p_34_1 = p_34_3 & p_2_1;
 assign g_34_1 = g_34_3 | (p_34_3 & g_2_1);
 assign p_34_2 = p_34_3 & p_2_2;
 assign g_34_2 = g_34_3 | (p_34_3 & g_2_2);
 assign p_34_3 = p_34_19 & p_18_3;
 assign g_34_3 = g_34_19 | (p_34_19 & g_18_3);
 assign p_34_4 = p_34_19 & p_18_4;
 assign g_34_4 = g_34_19 | (p_34_19 & g_18_4);
 assign p_34_5 = p_34_19 & p_18_5;
 assign g_34_5 = g_34_19 | (p_34_19 & g_18_5);
 assign p_34_6 = p_34_19 & p_18_6;
 assign g_34_6 = g_34_19 | (p_34_19 & g_18_6);
 assign p_34_7 = p_34_19 & p_18_7;
 assign g_34_7 = g_34_19 | (p_34_19 & g_18_7);
 assign p_34_8 = p_34_19 & p_18_8;
 assign g_34_8 = g_34_19 | (p_34_19 & g_18_8);
 assign p_34_9 = p_34_19 & p_18_9;
 assign g_34_9 = g_34_19 | (p_34_19 & g_18_9);
 assign p_34_10 = p_34_19 & p_18_10;
 assign g_34_10 = g_34_19 | (p_34_19 & g_18_10);
 assign p_34_11 = p_34_19 & p_18_11;
 assign g_34_11 = g_34_19 | (p_34_19 & g_18_11);
 assign p_34_12 = p_34_19 & p_18_12;
 assign g_34_12 = g_34_19 | (p_34_19 & g_18_12);
 assign p_34_13 = p_34_19 & p_18_13;
 assign g_34_13 = g_34_19 | (p_34_19 & g_18_13);
 assign p_34_14 = p_34_19 & p_18_14;
 assign g_34_14 = g_34_19 | (p_34_19 & g_18_14);
 assign p_34_15 = p_34_19 & p_18_15;
 assign g_34_15 = g_34_19 | (p_34_19 & g_18_15);
 assign p_34_16 = p_34_19 & p_18_16;
 assign g_34_16 = g_34_19 | (p_34_19 & g_18_16);
 assign p_34_17 = p_34_19 & p_18_17;
 assign g_34_17 = g_34_19 | (p_34_19 & g_18_17);
 assign p_34_18 = p_34_19 & p_18_18;
 assign g_34_18 = g_34_19 | (p_34_19 & g_18_18);
 assign p_34_19 = p_34_27 & p_26_19;
 assign g_34_19 = g_34_27 | (p_34_27 & g_26_19);
 assign p_34_20 = p_34_27 & p_26_20;
 assign g_34_20 = g_34_27 | (p_34_27 & g_26_20);
 assign p_34_21 = p_34_27 & p_26_21;
 assign g_34_21 = g_34_27 | (p_34_27 & g_26_21);
 assign p_34_22 = p_34_27 & p_26_22;
 assign g_34_22 = g_34_27 | (p_34_27 & g_26_22);
 assign p_34_23 = p_34_27 & p_26_23;
 assign g_34_23 = g_34_27 | (p_34_27 & g_26_23);
 assign p_34_24 = p_34_27 & p_26_24;
 assign g_34_24 = g_34_27 | (p_34_27 & g_26_24);
 assign p_34_25 = p_34_27 & p_26_25;
 assign g_34_25 = g_34_27 | (p_34_27 & g_26_25);
 assign p_34_26 = p_34_27 & p_26_26;
 assign g_34_26 = g_34_27 | (p_34_27 & g_26_26);
 assign p_34_27 = p_34_31 & p_30_27;
 assign g_34_27 = g_34_31 | (p_34_31 & g_30_27);
 assign p_34_28 = p_34_31 & p_30_28;
 assign g_34_28 = g_34_31 | (p_34_31 & g_30_28);
 assign p_34_29 = p_34_31 & p_30_29;
 assign g_34_29 = g_34_31 | (p_34_31 & g_30_29);
 assign p_34_30 = p_34_31 & p_30_30;
 assign g_34_30 = g_34_31 | (p_34_31 & g_30_30);
 assign p_34_31 = p_34_33 & p_32_31;
 assign g_34_31 = g_34_33 | (p_34_33 & g_32_31);
 assign p_34_32 = p_34_33 & p_32_32;
 assign g_34_32 = g_34_33 | (p_34_33 & g_32_32);
 assign p_34_33 = p_34_34 & p_33_33;
 assign g_34_33 = g_34_34 | (p_34_34 & g_33_33);
 assign sum[34] = p_34_34^ g_33_0;
 assign p_35_0 = p_35_4 & p_3_0;
 assign g_35_0 = g_35_4 | (p_35_4 & g_3_0);
 assign p_35_1 = p_35_4 & p_3_1;
 assign g_35_1 = g_35_4 | (p_35_4 & g_3_1);
 assign p_35_2 = p_35_4 & p_3_2;
 assign g_35_2 = g_35_4 | (p_35_4 & g_3_2);
 assign p_35_3 = p_35_4 & p_3_3;
 assign g_35_3 = g_35_4 | (p_35_4 & g_3_3);
 assign p_35_4 = p_35_20 & p_19_4;
 assign g_35_4 = g_35_20 | (p_35_20 & g_19_4);
 assign p_35_5 = p_35_20 & p_19_5;
 assign g_35_5 = g_35_20 | (p_35_20 & g_19_5);
 assign p_35_6 = p_35_20 & p_19_6;
 assign g_35_6 = g_35_20 | (p_35_20 & g_19_6);
 assign p_35_7 = p_35_20 & p_19_7;
 assign g_35_7 = g_35_20 | (p_35_20 & g_19_7);
 assign p_35_8 = p_35_20 & p_19_8;
 assign g_35_8 = g_35_20 | (p_35_20 & g_19_8);
 assign p_35_9 = p_35_20 & p_19_9;
 assign g_35_9 = g_35_20 | (p_35_20 & g_19_9);
 assign p_35_10 = p_35_20 & p_19_10;
 assign g_35_10 = g_35_20 | (p_35_20 & g_19_10);
 assign p_35_11 = p_35_20 & p_19_11;
 assign g_35_11 = g_35_20 | (p_35_20 & g_19_11);
 assign p_35_12 = p_35_20 & p_19_12;
 assign g_35_12 = g_35_20 | (p_35_20 & g_19_12);
 assign p_35_13 = p_35_20 & p_19_13;
 assign g_35_13 = g_35_20 | (p_35_20 & g_19_13);
 assign p_35_14 = p_35_20 & p_19_14;
 assign g_35_14 = g_35_20 | (p_35_20 & g_19_14);
 assign p_35_15 = p_35_20 & p_19_15;
 assign g_35_15 = g_35_20 | (p_35_20 & g_19_15);
 assign p_35_16 = p_35_20 & p_19_16;
 assign g_35_16 = g_35_20 | (p_35_20 & g_19_16);
 assign p_35_17 = p_35_20 & p_19_17;
 assign g_35_17 = g_35_20 | (p_35_20 & g_19_17);
 assign p_35_18 = p_35_20 & p_19_18;
 assign g_35_18 = g_35_20 | (p_35_20 & g_19_18);
 assign p_35_19 = p_35_20 & p_19_19;
 assign g_35_19 = g_35_20 | (p_35_20 & g_19_19);
 assign p_35_20 = p_35_28 & p_27_20;
 assign g_35_20 = g_35_28 | (p_35_28 & g_27_20);
 assign p_35_21 = p_35_28 & p_27_21;
 assign g_35_21 = g_35_28 | (p_35_28 & g_27_21);
 assign p_35_22 = p_35_28 & p_27_22;
 assign g_35_22 = g_35_28 | (p_35_28 & g_27_22);
 assign p_35_23 = p_35_28 & p_27_23;
 assign g_35_23 = g_35_28 | (p_35_28 & g_27_23);
 assign p_35_24 = p_35_28 & p_27_24;
 assign g_35_24 = g_35_28 | (p_35_28 & g_27_24);
 assign p_35_25 = p_35_28 & p_27_25;
 assign g_35_25 = g_35_28 | (p_35_28 & g_27_25);
 assign p_35_26 = p_35_28 & p_27_26;
 assign g_35_26 = g_35_28 | (p_35_28 & g_27_26);
 assign p_35_27 = p_35_28 & p_27_27;
 assign g_35_27 = g_35_28 | (p_35_28 & g_27_27);
 assign p_35_28 = p_35_32 & p_31_28;
 assign g_35_28 = g_35_32 | (p_35_32 & g_31_28);
 assign p_35_29 = p_35_32 & p_31_29;
 assign g_35_29 = g_35_32 | (p_35_32 & g_31_29);
 assign p_35_30 = p_35_32 & p_31_30;
 assign g_35_30 = g_35_32 | (p_35_32 & g_31_30);
 assign p_35_31 = p_35_32 & p_31_31;
 assign g_35_31 = g_35_32 | (p_35_32 & g_31_31);
 assign p_35_32 = p_35_34 & p_33_32;
 assign g_35_32 = g_35_34 | (p_35_34 & g_33_32);
 assign p_35_33 = p_35_34 & p_33_33;
 assign g_35_33 = g_35_34 | (p_35_34 & g_33_33);
 assign p_35_34 = p_35_35 & p_34_34;
 assign g_35_34 = g_35_35 | (p_35_35 & g_34_34);
 assign sum[35] = p_35_35^ g_34_0;
 assign p_36_0 = p_36_5 & p_4_0;
 assign g_36_0 = g_36_5 | (p_36_5 & g_4_0);
 assign p_36_1 = p_36_5 & p_4_1;
 assign g_36_1 = g_36_5 | (p_36_5 & g_4_1);
 assign p_36_2 = p_36_5 & p_4_2;
 assign g_36_2 = g_36_5 | (p_36_5 & g_4_2);
 assign p_36_3 = p_36_5 & p_4_3;
 assign g_36_3 = g_36_5 | (p_36_5 & g_4_3);
 assign p_36_4 = p_36_5 & p_4_4;
 assign g_36_4 = g_36_5 | (p_36_5 & g_4_4);
 assign p_36_5 = p_36_21 & p_20_5;
 assign g_36_5 = g_36_21 | (p_36_21 & g_20_5);
 assign p_36_6 = p_36_21 & p_20_6;
 assign g_36_6 = g_36_21 | (p_36_21 & g_20_6);
 assign p_36_7 = p_36_21 & p_20_7;
 assign g_36_7 = g_36_21 | (p_36_21 & g_20_7);
 assign p_36_8 = p_36_21 & p_20_8;
 assign g_36_8 = g_36_21 | (p_36_21 & g_20_8);
 assign p_36_9 = p_36_21 & p_20_9;
 assign g_36_9 = g_36_21 | (p_36_21 & g_20_9);
 assign p_36_10 = p_36_21 & p_20_10;
 assign g_36_10 = g_36_21 | (p_36_21 & g_20_10);
 assign p_36_11 = p_36_21 & p_20_11;
 assign g_36_11 = g_36_21 | (p_36_21 & g_20_11);
 assign p_36_12 = p_36_21 & p_20_12;
 assign g_36_12 = g_36_21 | (p_36_21 & g_20_12);
 assign p_36_13 = p_36_21 & p_20_13;
 assign g_36_13 = g_36_21 | (p_36_21 & g_20_13);
 assign p_36_14 = p_36_21 & p_20_14;
 assign g_36_14 = g_36_21 | (p_36_21 & g_20_14);
 assign p_36_15 = p_36_21 & p_20_15;
 assign g_36_15 = g_36_21 | (p_36_21 & g_20_15);
 assign p_36_16 = p_36_21 & p_20_16;
 assign g_36_16 = g_36_21 | (p_36_21 & g_20_16);
 assign p_36_17 = p_36_21 & p_20_17;
 assign g_36_17 = g_36_21 | (p_36_21 & g_20_17);
 assign p_36_18 = p_36_21 & p_20_18;
 assign g_36_18 = g_36_21 | (p_36_21 & g_20_18);
 assign p_36_19 = p_36_21 & p_20_19;
 assign g_36_19 = g_36_21 | (p_36_21 & g_20_19);
 assign p_36_20 = p_36_21 & p_20_20;
 assign g_36_20 = g_36_21 | (p_36_21 & g_20_20);
 assign p_36_21 = p_36_29 & p_28_21;
 assign g_36_21 = g_36_29 | (p_36_29 & g_28_21);
 assign p_36_22 = p_36_29 & p_28_22;
 assign g_36_22 = g_36_29 | (p_36_29 & g_28_22);
 assign p_36_23 = p_36_29 & p_28_23;
 assign g_36_23 = g_36_29 | (p_36_29 & g_28_23);
 assign p_36_24 = p_36_29 & p_28_24;
 assign g_36_24 = g_36_29 | (p_36_29 & g_28_24);
 assign p_36_25 = p_36_29 & p_28_25;
 assign g_36_25 = g_36_29 | (p_36_29 & g_28_25);
 assign p_36_26 = p_36_29 & p_28_26;
 assign g_36_26 = g_36_29 | (p_36_29 & g_28_26);
 assign p_36_27 = p_36_29 & p_28_27;
 assign g_36_27 = g_36_29 | (p_36_29 & g_28_27);
 assign p_36_28 = p_36_29 & p_28_28;
 assign g_36_28 = g_36_29 | (p_36_29 & g_28_28);
 assign p_36_29 = p_36_33 & p_32_29;
 assign g_36_29 = g_36_33 | (p_36_33 & g_32_29);
 assign p_36_30 = p_36_33 & p_32_30;
 assign g_36_30 = g_36_33 | (p_36_33 & g_32_30);
 assign p_36_31 = p_36_33 & p_32_31;
 assign g_36_31 = g_36_33 | (p_36_33 & g_32_31);
 assign p_36_32 = p_36_33 & p_32_32;
 assign g_36_32 = g_36_33 | (p_36_33 & g_32_32);
 assign p_36_33 = p_36_35 & p_34_33;
 assign g_36_33 = g_36_35 | (p_36_35 & g_34_33);
 assign p_36_34 = p_36_35 & p_34_34;
 assign g_36_34 = g_36_35 | (p_36_35 & g_34_34);
 assign p_36_35 = p_36_36 & p_35_35;
 assign g_36_35 = g_36_36 | (p_36_36 & g_35_35);
 assign sum[36] = p_36_36^ g_35_0;
 assign p_37_0 = p_37_6 & p_5_0;
 assign g_37_0 = g_37_6 | (p_37_6 & g_5_0);
 assign p_37_1 = p_37_6 & p_5_1;
 assign g_37_1 = g_37_6 | (p_37_6 & g_5_1);
 assign p_37_2 = p_37_6 & p_5_2;
 assign g_37_2 = g_37_6 | (p_37_6 & g_5_2);
 assign p_37_3 = p_37_6 & p_5_3;
 assign g_37_3 = g_37_6 | (p_37_6 & g_5_3);
 assign p_37_4 = p_37_6 & p_5_4;
 assign g_37_4 = g_37_6 | (p_37_6 & g_5_4);
 assign p_37_5 = p_37_6 & p_5_5;
 assign g_37_5 = g_37_6 | (p_37_6 & g_5_5);
 assign p_37_6 = p_37_22 & p_21_6;
 assign g_37_6 = g_37_22 | (p_37_22 & g_21_6);
 assign p_37_7 = p_37_22 & p_21_7;
 assign g_37_7 = g_37_22 | (p_37_22 & g_21_7);
 assign p_37_8 = p_37_22 & p_21_8;
 assign g_37_8 = g_37_22 | (p_37_22 & g_21_8);
 assign p_37_9 = p_37_22 & p_21_9;
 assign g_37_9 = g_37_22 | (p_37_22 & g_21_9);
 assign p_37_10 = p_37_22 & p_21_10;
 assign g_37_10 = g_37_22 | (p_37_22 & g_21_10);
 assign p_37_11 = p_37_22 & p_21_11;
 assign g_37_11 = g_37_22 | (p_37_22 & g_21_11);
 assign p_37_12 = p_37_22 & p_21_12;
 assign g_37_12 = g_37_22 | (p_37_22 & g_21_12);
 assign p_37_13 = p_37_22 & p_21_13;
 assign g_37_13 = g_37_22 | (p_37_22 & g_21_13);
 assign p_37_14 = p_37_22 & p_21_14;
 assign g_37_14 = g_37_22 | (p_37_22 & g_21_14);
 assign p_37_15 = p_37_22 & p_21_15;
 assign g_37_15 = g_37_22 | (p_37_22 & g_21_15);
 assign p_37_16 = p_37_22 & p_21_16;
 assign g_37_16 = g_37_22 | (p_37_22 & g_21_16);
 assign p_37_17 = p_37_22 & p_21_17;
 assign g_37_17 = g_37_22 | (p_37_22 & g_21_17);
 assign p_37_18 = p_37_22 & p_21_18;
 assign g_37_18 = g_37_22 | (p_37_22 & g_21_18);
 assign p_37_19 = p_37_22 & p_21_19;
 assign g_37_19 = g_37_22 | (p_37_22 & g_21_19);
 assign p_37_20 = p_37_22 & p_21_20;
 assign g_37_20 = g_37_22 | (p_37_22 & g_21_20);
 assign p_37_21 = p_37_22 & p_21_21;
 assign g_37_21 = g_37_22 | (p_37_22 & g_21_21);
 assign p_37_22 = p_37_30 & p_29_22;
 assign g_37_22 = g_37_30 | (p_37_30 & g_29_22);
 assign p_37_23 = p_37_30 & p_29_23;
 assign g_37_23 = g_37_30 | (p_37_30 & g_29_23);
 assign p_37_24 = p_37_30 & p_29_24;
 assign g_37_24 = g_37_30 | (p_37_30 & g_29_24);
 assign p_37_25 = p_37_30 & p_29_25;
 assign g_37_25 = g_37_30 | (p_37_30 & g_29_25);
 assign p_37_26 = p_37_30 & p_29_26;
 assign g_37_26 = g_37_30 | (p_37_30 & g_29_26);
 assign p_37_27 = p_37_30 & p_29_27;
 assign g_37_27 = g_37_30 | (p_37_30 & g_29_27);
 assign p_37_28 = p_37_30 & p_29_28;
 assign g_37_28 = g_37_30 | (p_37_30 & g_29_28);
 assign p_37_29 = p_37_30 & p_29_29;
 assign g_37_29 = g_37_30 | (p_37_30 & g_29_29);
 assign p_37_30 = p_37_34 & p_33_30;
 assign g_37_30 = g_37_34 | (p_37_34 & g_33_30);
 assign p_37_31 = p_37_34 & p_33_31;
 assign g_37_31 = g_37_34 | (p_37_34 & g_33_31);
 assign p_37_32 = p_37_34 & p_33_32;
 assign g_37_32 = g_37_34 | (p_37_34 & g_33_32);
 assign p_37_33 = p_37_34 & p_33_33;
 assign g_37_33 = g_37_34 | (p_37_34 & g_33_33);
 assign p_37_34 = p_37_36 & p_35_34;
 assign g_37_34 = g_37_36 | (p_37_36 & g_35_34);
 assign p_37_35 = p_37_36 & p_35_35;
 assign g_37_35 = g_37_36 | (p_37_36 & g_35_35);
 assign p_37_36 = p_37_37 & p_36_36;
 assign g_37_36 = g_37_37 | (p_37_37 & g_36_36);
 assign sum[37] = p_37_37^ g_36_0;
 assign p_38_0 = p_38_7 & p_6_0;
 assign g_38_0 = g_38_7 | (p_38_7 & g_6_0);
 assign p_38_1 = p_38_7 & p_6_1;
 assign g_38_1 = g_38_7 | (p_38_7 & g_6_1);
 assign p_38_2 = p_38_7 & p_6_2;
 assign g_38_2 = g_38_7 | (p_38_7 & g_6_2);
 assign p_38_3 = p_38_7 & p_6_3;
 assign g_38_3 = g_38_7 | (p_38_7 & g_6_3);
 assign p_38_4 = p_38_7 & p_6_4;
 assign g_38_4 = g_38_7 | (p_38_7 & g_6_4);
 assign p_38_5 = p_38_7 & p_6_5;
 assign g_38_5 = g_38_7 | (p_38_7 & g_6_5);
 assign p_38_6 = p_38_7 & p_6_6;
 assign g_38_6 = g_38_7 | (p_38_7 & g_6_6);
 assign p_38_7 = p_38_23 & p_22_7;
 assign g_38_7 = g_38_23 | (p_38_23 & g_22_7);
 assign p_38_8 = p_38_23 & p_22_8;
 assign g_38_8 = g_38_23 | (p_38_23 & g_22_8);
 assign p_38_9 = p_38_23 & p_22_9;
 assign g_38_9 = g_38_23 | (p_38_23 & g_22_9);
 assign p_38_10 = p_38_23 & p_22_10;
 assign g_38_10 = g_38_23 | (p_38_23 & g_22_10);
 assign p_38_11 = p_38_23 & p_22_11;
 assign g_38_11 = g_38_23 | (p_38_23 & g_22_11);
 assign p_38_12 = p_38_23 & p_22_12;
 assign g_38_12 = g_38_23 | (p_38_23 & g_22_12);
 assign p_38_13 = p_38_23 & p_22_13;
 assign g_38_13 = g_38_23 | (p_38_23 & g_22_13);
 assign p_38_14 = p_38_23 & p_22_14;
 assign g_38_14 = g_38_23 | (p_38_23 & g_22_14);
 assign p_38_15 = p_38_23 & p_22_15;
 assign g_38_15 = g_38_23 | (p_38_23 & g_22_15);
 assign p_38_16 = p_38_23 & p_22_16;
 assign g_38_16 = g_38_23 | (p_38_23 & g_22_16);
 assign p_38_17 = p_38_23 & p_22_17;
 assign g_38_17 = g_38_23 | (p_38_23 & g_22_17);
 assign p_38_18 = p_38_23 & p_22_18;
 assign g_38_18 = g_38_23 | (p_38_23 & g_22_18);
 assign p_38_19 = p_38_23 & p_22_19;
 assign g_38_19 = g_38_23 | (p_38_23 & g_22_19);
 assign p_38_20 = p_38_23 & p_22_20;
 assign g_38_20 = g_38_23 | (p_38_23 & g_22_20);
 assign p_38_21 = p_38_23 & p_22_21;
 assign g_38_21 = g_38_23 | (p_38_23 & g_22_21);
 assign p_38_22 = p_38_23 & p_22_22;
 assign g_38_22 = g_38_23 | (p_38_23 & g_22_22);
 assign p_38_23 = p_38_31 & p_30_23;
 assign g_38_23 = g_38_31 | (p_38_31 & g_30_23);
 assign p_38_24 = p_38_31 & p_30_24;
 assign g_38_24 = g_38_31 | (p_38_31 & g_30_24);
 assign p_38_25 = p_38_31 & p_30_25;
 assign g_38_25 = g_38_31 | (p_38_31 & g_30_25);
 assign p_38_26 = p_38_31 & p_30_26;
 assign g_38_26 = g_38_31 | (p_38_31 & g_30_26);
 assign p_38_27 = p_38_31 & p_30_27;
 assign g_38_27 = g_38_31 | (p_38_31 & g_30_27);
 assign p_38_28 = p_38_31 & p_30_28;
 assign g_38_28 = g_38_31 | (p_38_31 & g_30_28);
 assign p_38_29 = p_38_31 & p_30_29;
 assign g_38_29 = g_38_31 | (p_38_31 & g_30_29);
 assign p_38_30 = p_38_31 & p_30_30;
 assign g_38_30 = g_38_31 | (p_38_31 & g_30_30);
 assign p_38_31 = p_38_35 & p_34_31;
 assign g_38_31 = g_38_35 | (p_38_35 & g_34_31);
 assign p_38_32 = p_38_35 & p_34_32;
 assign g_38_32 = g_38_35 | (p_38_35 & g_34_32);
 assign p_38_33 = p_38_35 & p_34_33;
 assign g_38_33 = g_38_35 | (p_38_35 & g_34_33);
 assign p_38_34 = p_38_35 & p_34_34;
 assign g_38_34 = g_38_35 | (p_38_35 & g_34_34);
 assign p_38_35 = p_38_37 & p_36_35;
 assign g_38_35 = g_38_37 | (p_38_37 & g_36_35);
 assign p_38_36 = p_38_37 & p_36_36;
 assign g_38_36 = g_38_37 | (p_38_37 & g_36_36);
 assign p_38_37 = p_38_38 & p_37_37;
 assign g_38_37 = g_38_38 | (p_38_38 & g_37_37);
 assign sum[38] = p_38_38^ g_37_0;
 assign p_39_0 = p_39_8 & p_7_0;
 assign g_39_0 = g_39_8 | (p_39_8 & g_7_0);
 assign p_39_1 = p_39_8 & p_7_1;
 assign g_39_1 = g_39_8 | (p_39_8 & g_7_1);
 assign p_39_2 = p_39_8 & p_7_2;
 assign g_39_2 = g_39_8 | (p_39_8 & g_7_2);
 assign p_39_3 = p_39_8 & p_7_3;
 assign g_39_3 = g_39_8 | (p_39_8 & g_7_3);
 assign p_39_4 = p_39_8 & p_7_4;
 assign g_39_4 = g_39_8 | (p_39_8 & g_7_4);
 assign p_39_5 = p_39_8 & p_7_5;
 assign g_39_5 = g_39_8 | (p_39_8 & g_7_5);
 assign p_39_6 = p_39_8 & p_7_6;
 assign g_39_6 = g_39_8 | (p_39_8 & g_7_6);
 assign p_39_7 = p_39_8 & p_7_7;
 assign g_39_7 = g_39_8 | (p_39_8 & g_7_7);
 assign p_39_8 = p_39_24 & p_23_8;
 assign g_39_8 = g_39_24 | (p_39_24 & g_23_8);
 assign p_39_9 = p_39_24 & p_23_9;
 assign g_39_9 = g_39_24 | (p_39_24 & g_23_9);
 assign p_39_10 = p_39_24 & p_23_10;
 assign g_39_10 = g_39_24 | (p_39_24 & g_23_10);
 assign p_39_11 = p_39_24 & p_23_11;
 assign g_39_11 = g_39_24 | (p_39_24 & g_23_11);
 assign p_39_12 = p_39_24 & p_23_12;
 assign g_39_12 = g_39_24 | (p_39_24 & g_23_12);
 assign p_39_13 = p_39_24 & p_23_13;
 assign g_39_13 = g_39_24 | (p_39_24 & g_23_13);
 assign p_39_14 = p_39_24 & p_23_14;
 assign g_39_14 = g_39_24 | (p_39_24 & g_23_14);
 assign p_39_15 = p_39_24 & p_23_15;
 assign g_39_15 = g_39_24 | (p_39_24 & g_23_15);
 assign p_39_16 = p_39_24 & p_23_16;
 assign g_39_16 = g_39_24 | (p_39_24 & g_23_16);
 assign p_39_17 = p_39_24 & p_23_17;
 assign g_39_17 = g_39_24 | (p_39_24 & g_23_17);
 assign p_39_18 = p_39_24 & p_23_18;
 assign g_39_18 = g_39_24 | (p_39_24 & g_23_18);
 assign p_39_19 = p_39_24 & p_23_19;
 assign g_39_19 = g_39_24 | (p_39_24 & g_23_19);
 assign p_39_20 = p_39_24 & p_23_20;
 assign g_39_20 = g_39_24 | (p_39_24 & g_23_20);
 assign p_39_21 = p_39_24 & p_23_21;
 assign g_39_21 = g_39_24 | (p_39_24 & g_23_21);
 assign p_39_22 = p_39_24 & p_23_22;
 assign g_39_22 = g_39_24 | (p_39_24 & g_23_22);
 assign p_39_23 = p_39_24 & p_23_23;
 assign g_39_23 = g_39_24 | (p_39_24 & g_23_23);
 assign p_39_24 = p_39_32 & p_31_24;
 assign g_39_24 = g_39_32 | (p_39_32 & g_31_24);
 assign p_39_25 = p_39_32 & p_31_25;
 assign g_39_25 = g_39_32 | (p_39_32 & g_31_25);
 assign p_39_26 = p_39_32 & p_31_26;
 assign g_39_26 = g_39_32 | (p_39_32 & g_31_26);
 assign p_39_27 = p_39_32 & p_31_27;
 assign g_39_27 = g_39_32 | (p_39_32 & g_31_27);
 assign p_39_28 = p_39_32 & p_31_28;
 assign g_39_28 = g_39_32 | (p_39_32 & g_31_28);
 assign p_39_29 = p_39_32 & p_31_29;
 assign g_39_29 = g_39_32 | (p_39_32 & g_31_29);
 assign p_39_30 = p_39_32 & p_31_30;
 assign g_39_30 = g_39_32 | (p_39_32 & g_31_30);
 assign p_39_31 = p_39_32 & p_31_31;
 assign g_39_31 = g_39_32 | (p_39_32 & g_31_31);
 assign p_39_32 = p_39_36 & p_35_32;
 assign g_39_32 = g_39_36 | (p_39_36 & g_35_32);
 assign p_39_33 = p_39_36 & p_35_33;
 assign g_39_33 = g_39_36 | (p_39_36 & g_35_33);
 assign p_39_34 = p_39_36 & p_35_34;
 assign g_39_34 = g_39_36 | (p_39_36 & g_35_34);
 assign p_39_35 = p_39_36 & p_35_35;
 assign g_39_35 = g_39_36 | (p_39_36 & g_35_35);
 assign p_39_36 = p_39_38 & p_37_36;
 assign g_39_36 = g_39_38 | (p_39_38 & g_37_36);
 assign p_39_37 = p_39_38 & p_37_37;
 assign g_39_37 = g_39_38 | (p_39_38 & g_37_37);
 assign p_39_38 = p_39_39 & p_38_38;
 assign g_39_38 = g_39_39 | (p_39_39 & g_38_38);
 assign sum[39] = p_39_39^ g_38_0;
 assign p_40_0 = p_40_9 & p_8_0;
 assign g_40_0 = g_40_9 | (p_40_9 & g_8_0);
 assign p_40_1 = p_40_9 & p_8_1;
 assign g_40_1 = g_40_9 | (p_40_9 & g_8_1);
 assign p_40_2 = p_40_9 & p_8_2;
 assign g_40_2 = g_40_9 | (p_40_9 & g_8_2);
 assign p_40_3 = p_40_9 & p_8_3;
 assign g_40_3 = g_40_9 | (p_40_9 & g_8_3);
 assign p_40_4 = p_40_9 & p_8_4;
 assign g_40_4 = g_40_9 | (p_40_9 & g_8_4);
 assign p_40_5 = p_40_9 & p_8_5;
 assign g_40_5 = g_40_9 | (p_40_9 & g_8_5);
 assign p_40_6 = p_40_9 & p_8_6;
 assign g_40_6 = g_40_9 | (p_40_9 & g_8_6);
 assign p_40_7 = p_40_9 & p_8_7;
 assign g_40_7 = g_40_9 | (p_40_9 & g_8_7);
 assign p_40_8 = p_40_9 & p_8_8;
 assign g_40_8 = g_40_9 | (p_40_9 & g_8_8);
 assign p_40_9 = p_40_25 & p_24_9;
 assign g_40_9 = g_40_25 | (p_40_25 & g_24_9);
 assign p_40_10 = p_40_25 & p_24_10;
 assign g_40_10 = g_40_25 | (p_40_25 & g_24_10);
 assign p_40_11 = p_40_25 & p_24_11;
 assign g_40_11 = g_40_25 | (p_40_25 & g_24_11);
 assign p_40_12 = p_40_25 & p_24_12;
 assign g_40_12 = g_40_25 | (p_40_25 & g_24_12);
 assign p_40_13 = p_40_25 & p_24_13;
 assign g_40_13 = g_40_25 | (p_40_25 & g_24_13);
 assign p_40_14 = p_40_25 & p_24_14;
 assign g_40_14 = g_40_25 | (p_40_25 & g_24_14);
 assign p_40_15 = p_40_25 & p_24_15;
 assign g_40_15 = g_40_25 | (p_40_25 & g_24_15);
 assign p_40_16 = p_40_25 & p_24_16;
 assign g_40_16 = g_40_25 | (p_40_25 & g_24_16);
 assign p_40_17 = p_40_25 & p_24_17;
 assign g_40_17 = g_40_25 | (p_40_25 & g_24_17);
 assign p_40_18 = p_40_25 & p_24_18;
 assign g_40_18 = g_40_25 | (p_40_25 & g_24_18);
 assign p_40_19 = p_40_25 & p_24_19;
 assign g_40_19 = g_40_25 | (p_40_25 & g_24_19);
 assign p_40_20 = p_40_25 & p_24_20;
 assign g_40_20 = g_40_25 | (p_40_25 & g_24_20);
 assign p_40_21 = p_40_25 & p_24_21;
 assign g_40_21 = g_40_25 | (p_40_25 & g_24_21);
 assign p_40_22 = p_40_25 & p_24_22;
 assign g_40_22 = g_40_25 | (p_40_25 & g_24_22);
 assign p_40_23 = p_40_25 & p_24_23;
 assign g_40_23 = g_40_25 | (p_40_25 & g_24_23);
 assign p_40_24 = p_40_25 & p_24_24;
 assign g_40_24 = g_40_25 | (p_40_25 & g_24_24);
 assign p_40_25 = p_40_33 & p_32_25;
 assign g_40_25 = g_40_33 | (p_40_33 & g_32_25);
 assign p_40_26 = p_40_33 & p_32_26;
 assign g_40_26 = g_40_33 | (p_40_33 & g_32_26);
 assign p_40_27 = p_40_33 & p_32_27;
 assign g_40_27 = g_40_33 | (p_40_33 & g_32_27);
 assign p_40_28 = p_40_33 & p_32_28;
 assign g_40_28 = g_40_33 | (p_40_33 & g_32_28);
 assign p_40_29 = p_40_33 & p_32_29;
 assign g_40_29 = g_40_33 | (p_40_33 & g_32_29);
 assign p_40_30 = p_40_33 & p_32_30;
 assign g_40_30 = g_40_33 | (p_40_33 & g_32_30);
 assign p_40_31 = p_40_33 & p_32_31;
 assign g_40_31 = g_40_33 | (p_40_33 & g_32_31);
 assign p_40_32 = p_40_33 & p_32_32;
 assign g_40_32 = g_40_33 | (p_40_33 & g_32_32);
 assign p_40_33 = p_40_37 & p_36_33;
 assign g_40_33 = g_40_37 | (p_40_37 & g_36_33);
 assign p_40_34 = p_40_37 & p_36_34;
 assign g_40_34 = g_40_37 | (p_40_37 & g_36_34);
 assign p_40_35 = p_40_37 & p_36_35;
 assign g_40_35 = g_40_37 | (p_40_37 & g_36_35);
 assign p_40_36 = p_40_37 & p_36_36;
 assign g_40_36 = g_40_37 | (p_40_37 & g_36_36);
 assign p_40_37 = p_40_39 & p_38_37;
 assign g_40_37 = g_40_39 | (p_40_39 & g_38_37);
 assign p_40_38 = p_40_39 & p_38_38;
 assign g_40_38 = g_40_39 | (p_40_39 & g_38_38);
 assign p_40_39 = p_40_40 & p_39_39;
 assign g_40_39 = g_40_40 | (p_40_40 & g_39_39);
 assign sum[40] = p_40_40^ g_39_0;
 assign p_41_0 = p_41_10 & p_9_0;
 assign g_41_0 = g_41_10 | (p_41_10 & g_9_0);
 assign p_41_1 = p_41_10 & p_9_1;
 assign g_41_1 = g_41_10 | (p_41_10 & g_9_1);
 assign p_41_2 = p_41_10 & p_9_2;
 assign g_41_2 = g_41_10 | (p_41_10 & g_9_2);
 assign p_41_3 = p_41_10 & p_9_3;
 assign g_41_3 = g_41_10 | (p_41_10 & g_9_3);
 assign p_41_4 = p_41_10 & p_9_4;
 assign g_41_4 = g_41_10 | (p_41_10 & g_9_4);
 assign p_41_5 = p_41_10 & p_9_5;
 assign g_41_5 = g_41_10 | (p_41_10 & g_9_5);
 assign p_41_6 = p_41_10 & p_9_6;
 assign g_41_6 = g_41_10 | (p_41_10 & g_9_6);
 assign p_41_7 = p_41_10 & p_9_7;
 assign g_41_7 = g_41_10 | (p_41_10 & g_9_7);
 assign p_41_8 = p_41_10 & p_9_8;
 assign g_41_8 = g_41_10 | (p_41_10 & g_9_8);
 assign p_41_9 = p_41_10 & p_9_9;
 assign g_41_9 = g_41_10 | (p_41_10 & g_9_9);
 assign p_41_10 = p_41_26 & p_25_10;
 assign g_41_10 = g_41_26 | (p_41_26 & g_25_10);
 assign p_41_11 = p_41_26 & p_25_11;
 assign g_41_11 = g_41_26 | (p_41_26 & g_25_11);
 assign p_41_12 = p_41_26 & p_25_12;
 assign g_41_12 = g_41_26 | (p_41_26 & g_25_12);
 assign p_41_13 = p_41_26 & p_25_13;
 assign g_41_13 = g_41_26 | (p_41_26 & g_25_13);
 assign p_41_14 = p_41_26 & p_25_14;
 assign g_41_14 = g_41_26 | (p_41_26 & g_25_14);
 assign p_41_15 = p_41_26 & p_25_15;
 assign g_41_15 = g_41_26 | (p_41_26 & g_25_15);
 assign p_41_16 = p_41_26 & p_25_16;
 assign g_41_16 = g_41_26 | (p_41_26 & g_25_16);
 assign p_41_17 = p_41_26 & p_25_17;
 assign g_41_17 = g_41_26 | (p_41_26 & g_25_17);
 assign p_41_18 = p_41_26 & p_25_18;
 assign g_41_18 = g_41_26 | (p_41_26 & g_25_18);
 assign p_41_19 = p_41_26 & p_25_19;
 assign g_41_19 = g_41_26 | (p_41_26 & g_25_19);
 assign p_41_20 = p_41_26 & p_25_20;
 assign g_41_20 = g_41_26 | (p_41_26 & g_25_20);
 assign p_41_21 = p_41_26 & p_25_21;
 assign g_41_21 = g_41_26 | (p_41_26 & g_25_21);
 assign p_41_22 = p_41_26 & p_25_22;
 assign g_41_22 = g_41_26 | (p_41_26 & g_25_22);
 assign p_41_23 = p_41_26 & p_25_23;
 assign g_41_23 = g_41_26 | (p_41_26 & g_25_23);
 assign p_41_24 = p_41_26 & p_25_24;
 assign g_41_24 = g_41_26 | (p_41_26 & g_25_24);
 assign p_41_25 = p_41_26 & p_25_25;
 assign g_41_25 = g_41_26 | (p_41_26 & g_25_25);
 assign p_41_26 = p_41_34 & p_33_26;
 assign g_41_26 = g_41_34 | (p_41_34 & g_33_26);
 assign p_41_27 = p_41_34 & p_33_27;
 assign g_41_27 = g_41_34 | (p_41_34 & g_33_27);
 assign p_41_28 = p_41_34 & p_33_28;
 assign g_41_28 = g_41_34 | (p_41_34 & g_33_28);
 assign p_41_29 = p_41_34 & p_33_29;
 assign g_41_29 = g_41_34 | (p_41_34 & g_33_29);
 assign p_41_30 = p_41_34 & p_33_30;
 assign g_41_30 = g_41_34 | (p_41_34 & g_33_30);
 assign p_41_31 = p_41_34 & p_33_31;
 assign g_41_31 = g_41_34 | (p_41_34 & g_33_31);
 assign p_41_32 = p_41_34 & p_33_32;
 assign g_41_32 = g_41_34 | (p_41_34 & g_33_32);
 assign p_41_33 = p_41_34 & p_33_33;
 assign g_41_33 = g_41_34 | (p_41_34 & g_33_33);
 assign p_41_34 = p_41_38 & p_37_34;
 assign g_41_34 = g_41_38 | (p_41_38 & g_37_34);
 assign p_41_35 = p_41_38 & p_37_35;
 assign g_41_35 = g_41_38 | (p_41_38 & g_37_35);
 assign p_41_36 = p_41_38 & p_37_36;
 assign g_41_36 = g_41_38 | (p_41_38 & g_37_36);
 assign p_41_37 = p_41_38 & p_37_37;
 assign g_41_37 = g_41_38 | (p_41_38 & g_37_37);
 assign p_41_38 = p_41_40 & p_39_38;
 assign g_41_38 = g_41_40 | (p_41_40 & g_39_38);
 assign p_41_39 = p_41_40 & p_39_39;
 assign g_41_39 = g_41_40 | (p_41_40 & g_39_39);
 assign p_41_40 = p_41_41 & p_40_40;
 assign g_41_40 = g_41_41 | (p_41_41 & g_40_40);
 assign sum[41] = p_41_41^ g_40_0;
 assign p_42_0 = p_42_11 & p_10_0;
 assign g_42_0 = g_42_11 | (p_42_11 & g_10_0);
 assign p_42_1 = p_42_11 & p_10_1;
 assign g_42_1 = g_42_11 | (p_42_11 & g_10_1);
 assign p_42_2 = p_42_11 & p_10_2;
 assign g_42_2 = g_42_11 | (p_42_11 & g_10_2);
 assign p_42_3 = p_42_11 & p_10_3;
 assign g_42_3 = g_42_11 | (p_42_11 & g_10_3);
 assign p_42_4 = p_42_11 & p_10_4;
 assign g_42_4 = g_42_11 | (p_42_11 & g_10_4);
 assign p_42_5 = p_42_11 & p_10_5;
 assign g_42_5 = g_42_11 | (p_42_11 & g_10_5);
 assign p_42_6 = p_42_11 & p_10_6;
 assign g_42_6 = g_42_11 | (p_42_11 & g_10_6);
 assign p_42_7 = p_42_11 & p_10_7;
 assign g_42_7 = g_42_11 | (p_42_11 & g_10_7);
 assign p_42_8 = p_42_11 & p_10_8;
 assign g_42_8 = g_42_11 | (p_42_11 & g_10_8);
 assign p_42_9 = p_42_11 & p_10_9;
 assign g_42_9 = g_42_11 | (p_42_11 & g_10_9);
 assign p_42_10 = p_42_11 & p_10_10;
 assign g_42_10 = g_42_11 | (p_42_11 & g_10_10);
 assign p_42_11 = p_42_27 & p_26_11;
 assign g_42_11 = g_42_27 | (p_42_27 & g_26_11);
 assign p_42_12 = p_42_27 & p_26_12;
 assign g_42_12 = g_42_27 | (p_42_27 & g_26_12);
 assign p_42_13 = p_42_27 & p_26_13;
 assign g_42_13 = g_42_27 | (p_42_27 & g_26_13);
 assign p_42_14 = p_42_27 & p_26_14;
 assign g_42_14 = g_42_27 | (p_42_27 & g_26_14);
 assign p_42_15 = p_42_27 & p_26_15;
 assign g_42_15 = g_42_27 | (p_42_27 & g_26_15);
 assign p_42_16 = p_42_27 & p_26_16;
 assign g_42_16 = g_42_27 | (p_42_27 & g_26_16);
 assign p_42_17 = p_42_27 & p_26_17;
 assign g_42_17 = g_42_27 | (p_42_27 & g_26_17);
 assign p_42_18 = p_42_27 & p_26_18;
 assign g_42_18 = g_42_27 | (p_42_27 & g_26_18);
 assign p_42_19 = p_42_27 & p_26_19;
 assign g_42_19 = g_42_27 | (p_42_27 & g_26_19);
 assign p_42_20 = p_42_27 & p_26_20;
 assign g_42_20 = g_42_27 | (p_42_27 & g_26_20);
 assign p_42_21 = p_42_27 & p_26_21;
 assign g_42_21 = g_42_27 | (p_42_27 & g_26_21);
 assign p_42_22 = p_42_27 & p_26_22;
 assign g_42_22 = g_42_27 | (p_42_27 & g_26_22);
 assign p_42_23 = p_42_27 & p_26_23;
 assign g_42_23 = g_42_27 | (p_42_27 & g_26_23);
 assign p_42_24 = p_42_27 & p_26_24;
 assign g_42_24 = g_42_27 | (p_42_27 & g_26_24);
 assign p_42_25 = p_42_27 & p_26_25;
 assign g_42_25 = g_42_27 | (p_42_27 & g_26_25);
 assign p_42_26 = p_42_27 & p_26_26;
 assign g_42_26 = g_42_27 | (p_42_27 & g_26_26);
 assign p_42_27 = p_42_35 & p_34_27;
 assign g_42_27 = g_42_35 | (p_42_35 & g_34_27);
 assign p_42_28 = p_42_35 & p_34_28;
 assign g_42_28 = g_42_35 | (p_42_35 & g_34_28);
 assign p_42_29 = p_42_35 & p_34_29;
 assign g_42_29 = g_42_35 | (p_42_35 & g_34_29);
 assign p_42_30 = p_42_35 & p_34_30;
 assign g_42_30 = g_42_35 | (p_42_35 & g_34_30);
 assign p_42_31 = p_42_35 & p_34_31;
 assign g_42_31 = g_42_35 | (p_42_35 & g_34_31);
 assign p_42_32 = p_42_35 & p_34_32;
 assign g_42_32 = g_42_35 | (p_42_35 & g_34_32);
 assign p_42_33 = p_42_35 & p_34_33;
 assign g_42_33 = g_42_35 | (p_42_35 & g_34_33);
 assign p_42_34 = p_42_35 & p_34_34;
 assign g_42_34 = g_42_35 | (p_42_35 & g_34_34);
 assign p_42_35 = p_42_39 & p_38_35;
 assign g_42_35 = g_42_39 | (p_42_39 & g_38_35);
 assign p_42_36 = p_42_39 & p_38_36;
 assign g_42_36 = g_42_39 | (p_42_39 & g_38_36);
 assign p_42_37 = p_42_39 & p_38_37;
 assign g_42_37 = g_42_39 | (p_42_39 & g_38_37);
 assign p_42_38 = p_42_39 & p_38_38;
 assign g_42_38 = g_42_39 | (p_42_39 & g_38_38);
 assign p_42_39 = p_42_41 & p_40_39;
 assign g_42_39 = g_42_41 | (p_42_41 & g_40_39);
 assign p_42_40 = p_42_41 & p_40_40;
 assign g_42_40 = g_42_41 | (p_42_41 & g_40_40);
 assign p_42_41 = p_42_42 & p_41_41;
 assign g_42_41 = g_42_42 | (p_42_42 & g_41_41);
 assign sum[42] = p_42_42^ g_41_0;
 assign p_43_0 = p_43_12 & p_11_0;
 assign g_43_0 = g_43_12 | (p_43_12 & g_11_0);
 assign p_43_1 = p_43_12 & p_11_1;
 assign g_43_1 = g_43_12 | (p_43_12 & g_11_1);
 assign p_43_2 = p_43_12 & p_11_2;
 assign g_43_2 = g_43_12 | (p_43_12 & g_11_2);
 assign p_43_3 = p_43_12 & p_11_3;
 assign g_43_3 = g_43_12 | (p_43_12 & g_11_3);
 assign p_43_4 = p_43_12 & p_11_4;
 assign g_43_4 = g_43_12 | (p_43_12 & g_11_4);
 assign p_43_5 = p_43_12 & p_11_5;
 assign g_43_5 = g_43_12 | (p_43_12 & g_11_5);
 assign p_43_6 = p_43_12 & p_11_6;
 assign g_43_6 = g_43_12 | (p_43_12 & g_11_6);
 assign p_43_7 = p_43_12 & p_11_7;
 assign g_43_7 = g_43_12 | (p_43_12 & g_11_7);
 assign p_43_8 = p_43_12 & p_11_8;
 assign g_43_8 = g_43_12 | (p_43_12 & g_11_8);
 assign p_43_9 = p_43_12 & p_11_9;
 assign g_43_9 = g_43_12 | (p_43_12 & g_11_9);
 assign p_43_10 = p_43_12 & p_11_10;
 assign g_43_10 = g_43_12 | (p_43_12 & g_11_10);
 assign p_43_11 = p_43_12 & p_11_11;
 assign g_43_11 = g_43_12 | (p_43_12 & g_11_11);
 assign p_43_12 = p_43_28 & p_27_12;
 assign g_43_12 = g_43_28 | (p_43_28 & g_27_12);
 assign p_43_13 = p_43_28 & p_27_13;
 assign g_43_13 = g_43_28 | (p_43_28 & g_27_13);
 assign p_43_14 = p_43_28 & p_27_14;
 assign g_43_14 = g_43_28 | (p_43_28 & g_27_14);
 assign p_43_15 = p_43_28 & p_27_15;
 assign g_43_15 = g_43_28 | (p_43_28 & g_27_15);
 assign p_43_16 = p_43_28 & p_27_16;
 assign g_43_16 = g_43_28 | (p_43_28 & g_27_16);
 assign p_43_17 = p_43_28 & p_27_17;
 assign g_43_17 = g_43_28 | (p_43_28 & g_27_17);
 assign p_43_18 = p_43_28 & p_27_18;
 assign g_43_18 = g_43_28 | (p_43_28 & g_27_18);
 assign p_43_19 = p_43_28 & p_27_19;
 assign g_43_19 = g_43_28 | (p_43_28 & g_27_19);
 assign p_43_20 = p_43_28 & p_27_20;
 assign g_43_20 = g_43_28 | (p_43_28 & g_27_20);
 assign p_43_21 = p_43_28 & p_27_21;
 assign g_43_21 = g_43_28 | (p_43_28 & g_27_21);
 assign p_43_22 = p_43_28 & p_27_22;
 assign g_43_22 = g_43_28 | (p_43_28 & g_27_22);
 assign p_43_23 = p_43_28 & p_27_23;
 assign g_43_23 = g_43_28 | (p_43_28 & g_27_23);
 assign p_43_24 = p_43_28 & p_27_24;
 assign g_43_24 = g_43_28 | (p_43_28 & g_27_24);
 assign p_43_25 = p_43_28 & p_27_25;
 assign g_43_25 = g_43_28 | (p_43_28 & g_27_25);
 assign p_43_26 = p_43_28 & p_27_26;
 assign g_43_26 = g_43_28 | (p_43_28 & g_27_26);
 assign p_43_27 = p_43_28 & p_27_27;
 assign g_43_27 = g_43_28 | (p_43_28 & g_27_27);
 assign p_43_28 = p_43_36 & p_35_28;
 assign g_43_28 = g_43_36 | (p_43_36 & g_35_28);
 assign p_43_29 = p_43_36 & p_35_29;
 assign g_43_29 = g_43_36 | (p_43_36 & g_35_29);
 assign p_43_30 = p_43_36 & p_35_30;
 assign g_43_30 = g_43_36 | (p_43_36 & g_35_30);
 assign p_43_31 = p_43_36 & p_35_31;
 assign g_43_31 = g_43_36 | (p_43_36 & g_35_31);
 assign p_43_32 = p_43_36 & p_35_32;
 assign g_43_32 = g_43_36 | (p_43_36 & g_35_32);
 assign p_43_33 = p_43_36 & p_35_33;
 assign g_43_33 = g_43_36 | (p_43_36 & g_35_33);
 assign p_43_34 = p_43_36 & p_35_34;
 assign g_43_34 = g_43_36 | (p_43_36 & g_35_34);
 assign p_43_35 = p_43_36 & p_35_35;
 assign g_43_35 = g_43_36 | (p_43_36 & g_35_35);
 assign p_43_36 = p_43_40 & p_39_36;
 assign g_43_36 = g_43_40 | (p_43_40 & g_39_36);
 assign p_43_37 = p_43_40 & p_39_37;
 assign g_43_37 = g_43_40 | (p_43_40 & g_39_37);
 assign p_43_38 = p_43_40 & p_39_38;
 assign g_43_38 = g_43_40 | (p_43_40 & g_39_38);
 assign p_43_39 = p_43_40 & p_39_39;
 assign g_43_39 = g_43_40 | (p_43_40 & g_39_39);
 assign p_43_40 = p_43_42 & p_41_40;
 assign g_43_40 = g_43_42 | (p_43_42 & g_41_40);
 assign p_43_41 = p_43_42 & p_41_41;
 assign g_43_41 = g_43_42 | (p_43_42 & g_41_41);
 assign p_43_42 = p_43_43 & p_42_42;
 assign g_43_42 = g_43_43 | (p_43_43 & g_42_42);
 assign sum[43] = p_43_43^ g_42_0;
 assign p_44_0 = p_44_13 & p_12_0;
 assign g_44_0 = g_44_13 | (p_44_13 & g_12_0);
 assign p_44_1 = p_44_13 & p_12_1;
 assign g_44_1 = g_44_13 | (p_44_13 & g_12_1);
 assign p_44_2 = p_44_13 & p_12_2;
 assign g_44_2 = g_44_13 | (p_44_13 & g_12_2);
 assign p_44_3 = p_44_13 & p_12_3;
 assign g_44_3 = g_44_13 | (p_44_13 & g_12_3);
 assign p_44_4 = p_44_13 & p_12_4;
 assign g_44_4 = g_44_13 | (p_44_13 & g_12_4);
 assign p_44_5 = p_44_13 & p_12_5;
 assign g_44_5 = g_44_13 | (p_44_13 & g_12_5);
 assign p_44_6 = p_44_13 & p_12_6;
 assign g_44_6 = g_44_13 | (p_44_13 & g_12_6);
 assign p_44_7 = p_44_13 & p_12_7;
 assign g_44_7 = g_44_13 | (p_44_13 & g_12_7);
 assign p_44_8 = p_44_13 & p_12_8;
 assign g_44_8 = g_44_13 | (p_44_13 & g_12_8);
 assign p_44_9 = p_44_13 & p_12_9;
 assign g_44_9 = g_44_13 | (p_44_13 & g_12_9);
 assign p_44_10 = p_44_13 & p_12_10;
 assign g_44_10 = g_44_13 | (p_44_13 & g_12_10);
 assign p_44_11 = p_44_13 & p_12_11;
 assign g_44_11 = g_44_13 | (p_44_13 & g_12_11);
 assign p_44_12 = p_44_13 & p_12_12;
 assign g_44_12 = g_44_13 | (p_44_13 & g_12_12);
 assign p_44_13 = p_44_29 & p_28_13;
 assign g_44_13 = g_44_29 | (p_44_29 & g_28_13);
 assign p_44_14 = p_44_29 & p_28_14;
 assign g_44_14 = g_44_29 | (p_44_29 & g_28_14);
 assign p_44_15 = p_44_29 & p_28_15;
 assign g_44_15 = g_44_29 | (p_44_29 & g_28_15);
 assign p_44_16 = p_44_29 & p_28_16;
 assign g_44_16 = g_44_29 | (p_44_29 & g_28_16);
 assign p_44_17 = p_44_29 & p_28_17;
 assign g_44_17 = g_44_29 | (p_44_29 & g_28_17);
 assign p_44_18 = p_44_29 & p_28_18;
 assign g_44_18 = g_44_29 | (p_44_29 & g_28_18);
 assign p_44_19 = p_44_29 & p_28_19;
 assign g_44_19 = g_44_29 | (p_44_29 & g_28_19);
 assign p_44_20 = p_44_29 & p_28_20;
 assign g_44_20 = g_44_29 | (p_44_29 & g_28_20);
 assign p_44_21 = p_44_29 & p_28_21;
 assign g_44_21 = g_44_29 | (p_44_29 & g_28_21);
 assign p_44_22 = p_44_29 & p_28_22;
 assign g_44_22 = g_44_29 | (p_44_29 & g_28_22);
 assign p_44_23 = p_44_29 & p_28_23;
 assign g_44_23 = g_44_29 | (p_44_29 & g_28_23);
 assign p_44_24 = p_44_29 & p_28_24;
 assign g_44_24 = g_44_29 | (p_44_29 & g_28_24);
 assign p_44_25 = p_44_29 & p_28_25;
 assign g_44_25 = g_44_29 | (p_44_29 & g_28_25);
 assign p_44_26 = p_44_29 & p_28_26;
 assign g_44_26 = g_44_29 | (p_44_29 & g_28_26);
 assign p_44_27 = p_44_29 & p_28_27;
 assign g_44_27 = g_44_29 | (p_44_29 & g_28_27);
 assign p_44_28 = p_44_29 & p_28_28;
 assign g_44_28 = g_44_29 | (p_44_29 & g_28_28);
 assign p_44_29 = p_44_37 & p_36_29;
 assign g_44_29 = g_44_37 | (p_44_37 & g_36_29);
 assign p_44_30 = p_44_37 & p_36_30;
 assign g_44_30 = g_44_37 | (p_44_37 & g_36_30);
 assign p_44_31 = p_44_37 & p_36_31;
 assign g_44_31 = g_44_37 | (p_44_37 & g_36_31);
 assign p_44_32 = p_44_37 & p_36_32;
 assign g_44_32 = g_44_37 | (p_44_37 & g_36_32);
 assign p_44_33 = p_44_37 & p_36_33;
 assign g_44_33 = g_44_37 | (p_44_37 & g_36_33);
 assign p_44_34 = p_44_37 & p_36_34;
 assign g_44_34 = g_44_37 | (p_44_37 & g_36_34);
 assign p_44_35 = p_44_37 & p_36_35;
 assign g_44_35 = g_44_37 | (p_44_37 & g_36_35);
 assign p_44_36 = p_44_37 & p_36_36;
 assign g_44_36 = g_44_37 | (p_44_37 & g_36_36);
 assign p_44_37 = p_44_41 & p_40_37;
 assign g_44_37 = g_44_41 | (p_44_41 & g_40_37);
 assign p_44_38 = p_44_41 & p_40_38;
 assign g_44_38 = g_44_41 | (p_44_41 & g_40_38);
 assign p_44_39 = p_44_41 & p_40_39;
 assign g_44_39 = g_44_41 | (p_44_41 & g_40_39);
 assign p_44_40 = p_44_41 & p_40_40;
 assign g_44_40 = g_44_41 | (p_44_41 & g_40_40);
 assign p_44_41 = p_44_43 & p_42_41;
 assign g_44_41 = g_44_43 | (p_44_43 & g_42_41);
 assign p_44_42 = p_44_43 & p_42_42;
 assign g_44_42 = g_44_43 | (p_44_43 & g_42_42);
 assign p_44_43 = p_44_44 & p_43_43;
 assign g_44_43 = g_44_44 | (p_44_44 & g_43_43);
 assign sum[44] = p_44_44^ g_43_0;
 assign p_45_0 = p_45_14 & p_13_0;
 assign g_45_0 = g_45_14 | (p_45_14 & g_13_0);
 assign p_45_1 = p_45_14 & p_13_1;
 assign g_45_1 = g_45_14 | (p_45_14 & g_13_1);
 assign p_45_2 = p_45_14 & p_13_2;
 assign g_45_2 = g_45_14 | (p_45_14 & g_13_2);
 assign p_45_3 = p_45_14 & p_13_3;
 assign g_45_3 = g_45_14 | (p_45_14 & g_13_3);
 assign p_45_4 = p_45_14 & p_13_4;
 assign g_45_4 = g_45_14 | (p_45_14 & g_13_4);
 assign p_45_5 = p_45_14 & p_13_5;
 assign g_45_5 = g_45_14 | (p_45_14 & g_13_5);
 assign p_45_6 = p_45_14 & p_13_6;
 assign g_45_6 = g_45_14 | (p_45_14 & g_13_6);
 assign p_45_7 = p_45_14 & p_13_7;
 assign g_45_7 = g_45_14 | (p_45_14 & g_13_7);
 assign p_45_8 = p_45_14 & p_13_8;
 assign g_45_8 = g_45_14 | (p_45_14 & g_13_8);
 assign p_45_9 = p_45_14 & p_13_9;
 assign g_45_9 = g_45_14 | (p_45_14 & g_13_9);
 assign p_45_10 = p_45_14 & p_13_10;
 assign g_45_10 = g_45_14 | (p_45_14 & g_13_10);
 assign p_45_11 = p_45_14 & p_13_11;
 assign g_45_11 = g_45_14 | (p_45_14 & g_13_11);
 assign p_45_12 = p_45_14 & p_13_12;
 assign g_45_12 = g_45_14 | (p_45_14 & g_13_12);
 assign p_45_13 = p_45_14 & p_13_13;
 assign g_45_13 = g_45_14 | (p_45_14 & g_13_13);
 assign p_45_14 = p_45_30 & p_29_14;
 assign g_45_14 = g_45_30 | (p_45_30 & g_29_14);
 assign p_45_15 = p_45_30 & p_29_15;
 assign g_45_15 = g_45_30 | (p_45_30 & g_29_15);
 assign p_45_16 = p_45_30 & p_29_16;
 assign g_45_16 = g_45_30 | (p_45_30 & g_29_16);
 assign p_45_17 = p_45_30 & p_29_17;
 assign g_45_17 = g_45_30 | (p_45_30 & g_29_17);
 assign p_45_18 = p_45_30 & p_29_18;
 assign g_45_18 = g_45_30 | (p_45_30 & g_29_18);
 assign p_45_19 = p_45_30 & p_29_19;
 assign g_45_19 = g_45_30 | (p_45_30 & g_29_19);
 assign p_45_20 = p_45_30 & p_29_20;
 assign g_45_20 = g_45_30 | (p_45_30 & g_29_20);
 assign p_45_21 = p_45_30 & p_29_21;
 assign g_45_21 = g_45_30 | (p_45_30 & g_29_21);
 assign p_45_22 = p_45_30 & p_29_22;
 assign g_45_22 = g_45_30 | (p_45_30 & g_29_22);
 assign p_45_23 = p_45_30 & p_29_23;
 assign g_45_23 = g_45_30 | (p_45_30 & g_29_23);
 assign p_45_24 = p_45_30 & p_29_24;
 assign g_45_24 = g_45_30 | (p_45_30 & g_29_24);
 assign p_45_25 = p_45_30 & p_29_25;
 assign g_45_25 = g_45_30 | (p_45_30 & g_29_25);
 assign p_45_26 = p_45_30 & p_29_26;
 assign g_45_26 = g_45_30 | (p_45_30 & g_29_26);
 assign p_45_27 = p_45_30 & p_29_27;
 assign g_45_27 = g_45_30 | (p_45_30 & g_29_27);
 assign p_45_28 = p_45_30 & p_29_28;
 assign g_45_28 = g_45_30 | (p_45_30 & g_29_28);
 assign p_45_29 = p_45_30 & p_29_29;
 assign g_45_29 = g_45_30 | (p_45_30 & g_29_29);
 assign p_45_30 = p_45_38 & p_37_30;
 assign g_45_30 = g_45_38 | (p_45_38 & g_37_30);
 assign p_45_31 = p_45_38 & p_37_31;
 assign g_45_31 = g_45_38 | (p_45_38 & g_37_31);
 assign p_45_32 = p_45_38 & p_37_32;
 assign g_45_32 = g_45_38 | (p_45_38 & g_37_32);
 assign p_45_33 = p_45_38 & p_37_33;
 assign g_45_33 = g_45_38 | (p_45_38 & g_37_33);
 assign p_45_34 = p_45_38 & p_37_34;
 assign g_45_34 = g_45_38 | (p_45_38 & g_37_34);
 assign p_45_35 = p_45_38 & p_37_35;
 assign g_45_35 = g_45_38 | (p_45_38 & g_37_35);
 assign p_45_36 = p_45_38 & p_37_36;
 assign g_45_36 = g_45_38 | (p_45_38 & g_37_36);
 assign p_45_37 = p_45_38 & p_37_37;
 assign g_45_37 = g_45_38 | (p_45_38 & g_37_37);
 assign p_45_38 = p_45_42 & p_41_38;
 assign g_45_38 = g_45_42 | (p_45_42 & g_41_38);
 assign p_45_39 = p_45_42 & p_41_39;
 assign g_45_39 = g_45_42 | (p_45_42 & g_41_39);
 assign p_45_40 = p_45_42 & p_41_40;
 assign g_45_40 = g_45_42 | (p_45_42 & g_41_40);
 assign p_45_41 = p_45_42 & p_41_41;
 assign g_45_41 = g_45_42 | (p_45_42 & g_41_41);
 assign p_45_42 = p_45_44 & p_43_42;
 assign g_45_42 = g_45_44 | (p_45_44 & g_43_42);
 assign p_45_43 = p_45_44 & p_43_43;
 assign g_45_43 = g_45_44 | (p_45_44 & g_43_43);
 assign p_45_44 = p_45_45 & p_44_44;
 assign g_45_44 = g_45_45 | (p_45_45 & g_44_44);
 assign sum[45] = p_45_45^ g_44_0;
 assign p_46_0 = p_46_15 & p_14_0;
 assign g_46_0 = g_46_15 | (p_46_15 & g_14_0);
 assign p_46_1 = p_46_15 & p_14_1;
 assign g_46_1 = g_46_15 | (p_46_15 & g_14_1);
 assign p_46_2 = p_46_15 & p_14_2;
 assign g_46_2 = g_46_15 | (p_46_15 & g_14_2);
 assign p_46_3 = p_46_15 & p_14_3;
 assign g_46_3 = g_46_15 | (p_46_15 & g_14_3);
 assign p_46_4 = p_46_15 & p_14_4;
 assign g_46_4 = g_46_15 | (p_46_15 & g_14_4);
 assign p_46_5 = p_46_15 & p_14_5;
 assign g_46_5 = g_46_15 | (p_46_15 & g_14_5);
 assign p_46_6 = p_46_15 & p_14_6;
 assign g_46_6 = g_46_15 | (p_46_15 & g_14_6);
 assign p_46_7 = p_46_15 & p_14_7;
 assign g_46_7 = g_46_15 | (p_46_15 & g_14_7);
 assign p_46_8 = p_46_15 & p_14_8;
 assign g_46_8 = g_46_15 | (p_46_15 & g_14_8);
 assign p_46_9 = p_46_15 & p_14_9;
 assign g_46_9 = g_46_15 | (p_46_15 & g_14_9);
 assign p_46_10 = p_46_15 & p_14_10;
 assign g_46_10 = g_46_15 | (p_46_15 & g_14_10);
 assign p_46_11 = p_46_15 & p_14_11;
 assign g_46_11 = g_46_15 | (p_46_15 & g_14_11);
 assign p_46_12 = p_46_15 & p_14_12;
 assign g_46_12 = g_46_15 | (p_46_15 & g_14_12);
 assign p_46_13 = p_46_15 & p_14_13;
 assign g_46_13 = g_46_15 | (p_46_15 & g_14_13);
 assign p_46_14 = p_46_15 & p_14_14;
 assign g_46_14 = g_46_15 | (p_46_15 & g_14_14);
 assign p_46_15 = p_46_31 & p_30_15;
 assign g_46_15 = g_46_31 | (p_46_31 & g_30_15);
 assign p_46_16 = p_46_31 & p_30_16;
 assign g_46_16 = g_46_31 | (p_46_31 & g_30_16);
 assign p_46_17 = p_46_31 & p_30_17;
 assign g_46_17 = g_46_31 | (p_46_31 & g_30_17);
 assign p_46_18 = p_46_31 & p_30_18;
 assign g_46_18 = g_46_31 | (p_46_31 & g_30_18);
 assign p_46_19 = p_46_31 & p_30_19;
 assign g_46_19 = g_46_31 | (p_46_31 & g_30_19);
 assign p_46_20 = p_46_31 & p_30_20;
 assign g_46_20 = g_46_31 | (p_46_31 & g_30_20);
 assign p_46_21 = p_46_31 & p_30_21;
 assign g_46_21 = g_46_31 | (p_46_31 & g_30_21);
 assign p_46_22 = p_46_31 & p_30_22;
 assign g_46_22 = g_46_31 | (p_46_31 & g_30_22);
 assign p_46_23 = p_46_31 & p_30_23;
 assign g_46_23 = g_46_31 | (p_46_31 & g_30_23);
 assign p_46_24 = p_46_31 & p_30_24;
 assign g_46_24 = g_46_31 | (p_46_31 & g_30_24);
 assign p_46_25 = p_46_31 & p_30_25;
 assign g_46_25 = g_46_31 | (p_46_31 & g_30_25);
 assign p_46_26 = p_46_31 & p_30_26;
 assign g_46_26 = g_46_31 | (p_46_31 & g_30_26);
 assign p_46_27 = p_46_31 & p_30_27;
 assign g_46_27 = g_46_31 | (p_46_31 & g_30_27);
 assign p_46_28 = p_46_31 & p_30_28;
 assign g_46_28 = g_46_31 | (p_46_31 & g_30_28);
 assign p_46_29 = p_46_31 & p_30_29;
 assign g_46_29 = g_46_31 | (p_46_31 & g_30_29);
 assign p_46_30 = p_46_31 & p_30_30;
 assign g_46_30 = g_46_31 | (p_46_31 & g_30_30);
 assign p_46_31 = p_46_39 & p_38_31;
 assign g_46_31 = g_46_39 | (p_46_39 & g_38_31);
 assign p_46_32 = p_46_39 & p_38_32;
 assign g_46_32 = g_46_39 | (p_46_39 & g_38_32);
 assign p_46_33 = p_46_39 & p_38_33;
 assign g_46_33 = g_46_39 | (p_46_39 & g_38_33);
 assign p_46_34 = p_46_39 & p_38_34;
 assign g_46_34 = g_46_39 | (p_46_39 & g_38_34);
 assign p_46_35 = p_46_39 & p_38_35;
 assign g_46_35 = g_46_39 | (p_46_39 & g_38_35);
 assign p_46_36 = p_46_39 & p_38_36;
 assign g_46_36 = g_46_39 | (p_46_39 & g_38_36);
 assign p_46_37 = p_46_39 & p_38_37;
 assign g_46_37 = g_46_39 | (p_46_39 & g_38_37);
 assign p_46_38 = p_46_39 & p_38_38;
 assign g_46_38 = g_46_39 | (p_46_39 & g_38_38);
 assign p_46_39 = p_46_43 & p_42_39;
 assign g_46_39 = g_46_43 | (p_46_43 & g_42_39);
 assign p_46_40 = p_46_43 & p_42_40;
 assign g_46_40 = g_46_43 | (p_46_43 & g_42_40);
 assign p_46_41 = p_46_43 & p_42_41;
 assign g_46_41 = g_46_43 | (p_46_43 & g_42_41);
 assign p_46_42 = p_46_43 & p_42_42;
 assign g_46_42 = g_46_43 | (p_46_43 & g_42_42);
 assign p_46_43 = p_46_45 & p_44_43;
 assign g_46_43 = g_46_45 | (p_46_45 & g_44_43);
 assign p_46_44 = p_46_45 & p_44_44;
 assign g_46_44 = g_46_45 | (p_46_45 & g_44_44);
 assign p_46_45 = p_46_46 & p_45_45;
 assign g_46_45 = g_46_46 | (p_46_46 & g_45_45);
 assign sum[46] = p_46_46^ g_45_0;
 assign p_47_0 = p_47_16 & p_15_0;
 assign g_47_0 = g_47_16 | (p_47_16 & g_15_0);
 assign p_47_1 = p_47_16 & p_15_1;
 assign g_47_1 = g_47_16 | (p_47_16 & g_15_1);
 assign p_47_2 = p_47_16 & p_15_2;
 assign g_47_2 = g_47_16 | (p_47_16 & g_15_2);
 assign p_47_3 = p_47_16 & p_15_3;
 assign g_47_3 = g_47_16 | (p_47_16 & g_15_3);
 assign p_47_4 = p_47_16 & p_15_4;
 assign g_47_4 = g_47_16 | (p_47_16 & g_15_4);
 assign p_47_5 = p_47_16 & p_15_5;
 assign g_47_5 = g_47_16 | (p_47_16 & g_15_5);
 assign p_47_6 = p_47_16 & p_15_6;
 assign g_47_6 = g_47_16 | (p_47_16 & g_15_6);
 assign p_47_7 = p_47_16 & p_15_7;
 assign g_47_7 = g_47_16 | (p_47_16 & g_15_7);
 assign p_47_8 = p_47_16 & p_15_8;
 assign g_47_8 = g_47_16 | (p_47_16 & g_15_8);
 assign p_47_9 = p_47_16 & p_15_9;
 assign g_47_9 = g_47_16 | (p_47_16 & g_15_9);
 assign p_47_10 = p_47_16 & p_15_10;
 assign g_47_10 = g_47_16 | (p_47_16 & g_15_10);
 assign p_47_11 = p_47_16 & p_15_11;
 assign g_47_11 = g_47_16 | (p_47_16 & g_15_11);
 assign p_47_12 = p_47_16 & p_15_12;
 assign g_47_12 = g_47_16 | (p_47_16 & g_15_12);
 assign p_47_13 = p_47_16 & p_15_13;
 assign g_47_13 = g_47_16 | (p_47_16 & g_15_13);
 assign p_47_14 = p_47_16 & p_15_14;
 assign g_47_14 = g_47_16 | (p_47_16 & g_15_14);
 assign p_47_15 = p_47_16 & p_15_15;
 assign g_47_15 = g_47_16 | (p_47_16 & g_15_15);
 assign p_47_16 = p_47_32 & p_31_16;
 assign g_47_16 = g_47_32 | (p_47_32 & g_31_16);
 assign p_47_17 = p_47_32 & p_31_17;
 assign g_47_17 = g_47_32 | (p_47_32 & g_31_17);
 assign p_47_18 = p_47_32 & p_31_18;
 assign g_47_18 = g_47_32 | (p_47_32 & g_31_18);
 assign p_47_19 = p_47_32 & p_31_19;
 assign g_47_19 = g_47_32 | (p_47_32 & g_31_19);
 assign p_47_20 = p_47_32 & p_31_20;
 assign g_47_20 = g_47_32 | (p_47_32 & g_31_20);
 assign p_47_21 = p_47_32 & p_31_21;
 assign g_47_21 = g_47_32 | (p_47_32 & g_31_21);
 assign p_47_22 = p_47_32 & p_31_22;
 assign g_47_22 = g_47_32 | (p_47_32 & g_31_22);
 assign p_47_23 = p_47_32 & p_31_23;
 assign g_47_23 = g_47_32 | (p_47_32 & g_31_23);
 assign p_47_24 = p_47_32 & p_31_24;
 assign g_47_24 = g_47_32 | (p_47_32 & g_31_24);
 assign p_47_25 = p_47_32 & p_31_25;
 assign g_47_25 = g_47_32 | (p_47_32 & g_31_25);
 assign p_47_26 = p_47_32 & p_31_26;
 assign g_47_26 = g_47_32 | (p_47_32 & g_31_26);
 assign p_47_27 = p_47_32 & p_31_27;
 assign g_47_27 = g_47_32 | (p_47_32 & g_31_27);
 assign p_47_28 = p_47_32 & p_31_28;
 assign g_47_28 = g_47_32 | (p_47_32 & g_31_28);
 assign p_47_29 = p_47_32 & p_31_29;
 assign g_47_29 = g_47_32 | (p_47_32 & g_31_29);
 assign p_47_30 = p_47_32 & p_31_30;
 assign g_47_30 = g_47_32 | (p_47_32 & g_31_30);
 assign p_47_31 = p_47_32 & p_31_31;
 assign g_47_31 = g_47_32 | (p_47_32 & g_31_31);
 assign p_47_32 = p_47_40 & p_39_32;
 assign g_47_32 = g_47_40 | (p_47_40 & g_39_32);
 assign p_47_33 = p_47_40 & p_39_33;
 assign g_47_33 = g_47_40 | (p_47_40 & g_39_33);
 assign p_47_34 = p_47_40 & p_39_34;
 assign g_47_34 = g_47_40 | (p_47_40 & g_39_34);
 assign p_47_35 = p_47_40 & p_39_35;
 assign g_47_35 = g_47_40 | (p_47_40 & g_39_35);
 assign p_47_36 = p_47_40 & p_39_36;
 assign g_47_36 = g_47_40 | (p_47_40 & g_39_36);
 assign p_47_37 = p_47_40 & p_39_37;
 assign g_47_37 = g_47_40 | (p_47_40 & g_39_37);
 assign p_47_38 = p_47_40 & p_39_38;
 assign g_47_38 = g_47_40 | (p_47_40 & g_39_38);
 assign p_47_39 = p_47_40 & p_39_39;
 assign g_47_39 = g_47_40 | (p_47_40 & g_39_39);
 assign p_47_40 = p_47_44 & p_43_40;
 assign g_47_40 = g_47_44 | (p_47_44 & g_43_40);
 assign p_47_41 = p_47_44 & p_43_41;
 assign g_47_41 = g_47_44 | (p_47_44 & g_43_41);
 assign p_47_42 = p_47_44 & p_43_42;
 assign g_47_42 = g_47_44 | (p_47_44 & g_43_42);
 assign p_47_43 = p_47_44 & p_43_43;
 assign g_47_43 = g_47_44 | (p_47_44 & g_43_43);
 assign p_47_44 = p_47_46 & p_45_44;
 assign g_47_44 = g_47_46 | (p_47_46 & g_45_44);
 assign p_47_45 = p_47_46 & p_45_45;
 assign g_47_45 = g_47_46 | (p_47_46 & g_45_45);
 assign p_47_46 = p_47_47 & p_46_46;
 assign g_47_46 = g_47_47 | (p_47_47 & g_46_46);
 assign sum[47] = p_47_47^ g_46_0;
 assign p_48_0 = p_48_17 & p_16_0;
 assign g_48_0 = g_48_17 | (p_48_17 & g_16_0);
 assign p_48_1 = p_48_17 & p_16_1;
 assign g_48_1 = g_48_17 | (p_48_17 & g_16_1);
 assign p_48_2 = p_48_17 & p_16_2;
 assign g_48_2 = g_48_17 | (p_48_17 & g_16_2);
 assign p_48_3 = p_48_17 & p_16_3;
 assign g_48_3 = g_48_17 | (p_48_17 & g_16_3);
 assign p_48_4 = p_48_17 & p_16_4;
 assign g_48_4 = g_48_17 | (p_48_17 & g_16_4);
 assign p_48_5 = p_48_17 & p_16_5;
 assign g_48_5 = g_48_17 | (p_48_17 & g_16_5);
 assign p_48_6 = p_48_17 & p_16_6;
 assign g_48_6 = g_48_17 | (p_48_17 & g_16_6);
 assign p_48_7 = p_48_17 & p_16_7;
 assign g_48_7 = g_48_17 | (p_48_17 & g_16_7);
 assign p_48_8 = p_48_17 & p_16_8;
 assign g_48_8 = g_48_17 | (p_48_17 & g_16_8);
 assign p_48_9 = p_48_17 & p_16_9;
 assign g_48_9 = g_48_17 | (p_48_17 & g_16_9);
 assign p_48_10 = p_48_17 & p_16_10;
 assign g_48_10 = g_48_17 | (p_48_17 & g_16_10);
 assign p_48_11 = p_48_17 & p_16_11;
 assign g_48_11 = g_48_17 | (p_48_17 & g_16_11);
 assign p_48_12 = p_48_17 & p_16_12;
 assign g_48_12 = g_48_17 | (p_48_17 & g_16_12);
 assign p_48_13 = p_48_17 & p_16_13;
 assign g_48_13 = g_48_17 | (p_48_17 & g_16_13);
 assign p_48_14 = p_48_17 & p_16_14;
 assign g_48_14 = g_48_17 | (p_48_17 & g_16_14);
 assign p_48_15 = p_48_17 & p_16_15;
 assign g_48_15 = g_48_17 | (p_48_17 & g_16_15);
 assign p_48_16 = p_48_17 & p_16_16;
 assign g_48_16 = g_48_17 | (p_48_17 & g_16_16);
 assign p_48_17 = p_48_33 & p_32_17;
 assign g_48_17 = g_48_33 | (p_48_33 & g_32_17);
 assign p_48_18 = p_48_33 & p_32_18;
 assign g_48_18 = g_48_33 | (p_48_33 & g_32_18);
 assign p_48_19 = p_48_33 & p_32_19;
 assign g_48_19 = g_48_33 | (p_48_33 & g_32_19);
 assign p_48_20 = p_48_33 & p_32_20;
 assign g_48_20 = g_48_33 | (p_48_33 & g_32_20);
 assign p_48_21 = p_48_33 & p_32_21;
 assign g_48_21 = g_48_33 | (p_48_33 & g_32_21);
 assign p_48_22 = p_48_33 & p_32_22;
 assign g_48_22 = g_48_33 | (p_48_33 & g_32_22);
 assign p_48_23 = p_48_33 & p_32_23;
 assign g_48_23 = g_48_33 | (p_48_33 & g_32_23);
 assign p_48_24 = p_48_33 & p_32_24;
 assign g_48_24 = g_48_33 | (p_48_33 & g_32_24);
 assign p_48_25 = p_48_33 & p_32_25;
 assign g_48_25 = g_48_33 | (p_48_33 & g_32_25);
 assign p_48_26 = p_48_33 & p_32_26;
 assign g_48_26 = g_48_33 | (p_48_33 & g_32_26);
 assign p_48_27 = p_48_33 & p_32_27;
 assign g_48_27 = g_48_33 | (p_48_33 & g_32_27);
 assign p_48_28 = p_48_33 & p_32_28;
 assign g_48_28 = g_48_33 | (p_48_33 & g_32_28);
 assign p_48_29 = p_48_33 & p_32_29;
 assign g_48_29 = g_48_33 | (p_48_33 & g_32_29);
 assign p_48_30 = p_48_33 & p_32_30;
 assign g_48_30 = g_48_33 | (p_48_33 & g_32_30);
 assign p_48_31 = p_48_33 & p_32_31;
 assign g_48_31 = g_48_33 | (p_48_33 & g_32_31);
 assign p_48_32 = p_48_33 & p_32_32;
 assign g_48_32 = g_48_33 | (p_48_33 & g_32_32);
 assign p_48_33 = p_48_41 & p_40_33;
 assign g_48_33 = g_48_41 | (p_48_41 & g_40_33);
 assign p_48_34 = p_48_41 & p_40_34;
 assign g_48_34 = g_48_41 | (p_48_41 & g_40_34);
 assign p_48_35 = p_48_41 & p_40_35;
 assign g_48_35 = g_48_41 | (p_48_41 & g_40_35);
 assign p_48_36 = p_48_41 & p_40_36;
 assign g_48_36 = g_48_41 | (p_48_41 & g_40_36);
 assign p_48_37 = p_48_41 & p_40_37;
 assign g_48_37 = g_48_41 | (p_48_41 & g_40_37);
 assign p_48_38 = p_48_41 & p_40_38;
 assign g_48_38 = g_48_41 | (p_48_41 & g_40_38);
 assign p_48_39 = p_48_41 & p_40_39;
 assign g_48_39 = g_48_41 | (p_48_41 & g_40_39);
 assign p_48_40 = p_48_41 & p_40_40;
 assign g_48_40 = g_48_41 | (p_48_41 & g_40_40);
 assign p_48_41 = p_48_45 & p_44_41;
 assign g_48_41 = g_48_45 | (p_48_45 & g_44_41);
 assign p_48_42 = p_48_45 & p_44_42;
 assign g_48_42 = g_48_45 | (p_48_45 & g_44_42);
 assign p_48_43 = p_48_45 & p_44_43;
 assign g_48_43 = g_48_45 | (p_48_45 & g_44_43);
 assign p_48_44 = p_48_45 & p_44_44;
 assign g_48_44 = g_48_45 | (p_48_45 & g_44_44);
 assign p_48_45 = p_48_47 & p_46_45;
 assign g_48_45 = g_48_47 | (p_48_47 & g_46_45);
 assign p_48_46 = p_48_47 & p_46_46;
 assign g_48_46 = g_48_47 | (p_48_47 & g_46_46);
 assign p_48_47 = p_48_48 & p_47_47;
 assign g_48_47 = g_48_48 | (p_48_48 & g_47_47);
 assign sum[48] = p_48_48^ g_47_0;
 assign p_49_0 = p_49_18 & p_17_0;
 assign g_49_0 = g_49_18 | (p_49_18 & g_17_0);
 assign p_49_1 = p_49_18 & p_17_1;
 assign g_49_1 = g_49_18 | (p_49_18 & g_17_1);
 assign p_49_2 = p_49_18 & p_17_2;
 assign g_49_2 = g_49_18 | (p_49_18 & g_17_2);
 assign p_49_3 = p_49_18 & p_17_3;
 assign g_49_3 = g_49_18 | (p_49_18 & g_17_3);
 assign p_49_4 = p_49_18 & p_17_4;
 assign g_49_4 = g_49_18 | (p_49_18 & g_17_4);
 assign p_49_5 = p_49_18 & p_17_5;
 assign g_49_5 = g_49_18 | (p_49_18 & g_17_5);
 assign p_49_6 = p_49_18 & p_17_6;
 assign g_49_6 = g_49_18 | (p_49_18 & g_17_6);
 assign p_49_7 = p_49_18 & p_17_7;
 assign g_49_7 = g_49_18 | (p_49_18 & g_17_7);
 assign p_49_8 = p_49_18 & p_17_8;
 assign g_49_8 = g_49_18 | (p_49_18 & g_17_8);
 assign p_49_9 = p_49_18 & p_17_9;
 assign g_49_9 = g_49_18 | (p_49_18 & g_17_9);
 assign p_49_10 = p_49_18 & p_17_10;
 assign g_49_10 = g_49_18 | (p_49_18 & g_17_10);
 assign p_49_11 = p_49_18 & p_17_11;
 assign g_49_11 = g_49_18 | (p_49_18 & g_17_11);
 assign p_49_12 = p_49_18 & p_17_12;
 assign g_49_12 = g_49_18 | (p_49_18 & g_17_12);
 assign p_49_13 = p_49_18 & p_17_13;
 assign g_49_13 = g_49_18 | (p_49_18 & g_17_13);
 assign p_49_14 = p_49_18 & p_17_14;
 assign g_49_14 = g_49_18 | (p_49_18 & g_17_14);
 assign p_49_15 = p_49_18 & p_17_15;
 assign g_49_15 = g_49_18 | (p_49_18 & g_17_15);
 assign p_49_16 = p_49_18 & p_17_16;
 assign g_49_16 = g_49_18 | (p_49_18 & g_17_16);
 assign p_49_17 = p_49_18 & p_17_17;
 assign g_49_17 = g_49_18 | (p_49_18 & g_17_17);
 assign p_49_18 = p_49_34 & p_33_18;
 assign g_49_18 = g_49_34 | (p_49_34 & g_33_18);
 assign p_49_19 = p_49_34 & p_33_19;
 assign g_49_19 = g_49_34 | (p_49_34 & g_33_19);
 assign p_49_20 = p_49_34 & p_33_20;
 assign g_49_20 = g_49_34 | (p_49_34 & g_33_20);
 assign p_49_21 = p_49_34 & p_33_21;
 assign g_49_21 = g_49_34 | (p_49_34 & g_33_21);
 assign p_49_22 = p_49_34 & p_33_22;
 assign g_49_22 = g_49_34 | (p_49_34 & g_33_22);
 assign p_49_23 = p_49_34 & p_33_23;
 assign g_49_23 = g_49_34 | (p_49_34 & g_33_23);
 assign p_49_24 = p_49_34 & p_33_24;
 assign g_49_24 = g_49_34 | (p_49_34 & g_33_24);
 assign p_49_25 = p_49_34 & p_33_25;
 assign g_49_25 = g_49_34 | (p_49_34 & g_33_25);
 assign p_49_26 = p_49_34 & p_33_26;
 assign g_49_26 = g_49_34 | (p_49_34 & g_33_26);
 assign p_49_27 = p_49_34 & p_33_27;
 assign g_49_27 = g_49_34 | (p_49_34 & g_33_27);
 assign p_49_28 = p_49_34 & p_33_28;
 assign g_49_28 = g_49_34 | (p_49_34 & g_33_28);
 assign p_49_29 = p_49_34 & p_33_29;
 assign g_49_29 = g_49_34 | (p_49_34 & g_33_29);
 assign p_49_30 = p_49_34 & p_33_30;
 assign g_49_30 = g_49_34 | (p_49_34 & g_33_30);
 assign p_49_31 = p_49_34 & p_33_31;
 assign g_49_31 = g_49_34 | (p_49_34 & g_33_31);
 assign p_49_32 = p_49_34 & p_33_32;
 assign g_49_32 = g_49_34 | (p_49_34 & g_33_32);
 assign p_49_33 = p_49_34 & p_33_33;
 assign g_49_33 = g_49_34 | (p_49_34 & g_33_33);
 assign p_49_34 = p_49_42 & p_41_34;
 assign g_49_34 = g_49_42 | (p_49_42 & g_41_34);
 assign p_49_35 = p_49_42 & p_41_35;
 assign g_49_35 = g_49_42 | (p_49_42 & g_41_35);
 assign p_49_36 = p_49_42 & p_41_36;
 assign g_49_36 = g_49_42 | (p_49_42 & g_41_36);
 assign p_49_37 = p_49_42 & p_41_37;
 assign g_49_37 = g_49_42 | (p_49_42 & g_41_37);
 assign p_49_38 = p_49_42 & p_41_38;
 assign g_49_38 = g_49_42 | (p_49_42 & g_41_38);
 assign p_49_39 = p_49_42 & p_41_39;
 assign g_49_39 = g_49_42 | (p_49_42 & g_41_39);
 assign p_49_40 = p_49_42 & p_41_40;
 assign g_49_40 = g_49_42 | (p_49_42 & g_41_40);
 assign p_49_41 = p_49_42 & p_41_41;
 assign g_49_41 = g_49_42 | (p_49_42 & g_41_41);
 assign p_49_42 = p_49_46 & p_45_42;
 assign g_49_42 = g_49_46 | (p_49_46 & g_45_42);
 assign p_49_43 = p_49_46 & p_45_43;
 assign g_49_43 = g_49_46 | (p_49_46 & g_45_43);
 assign p_49_44 = p_49_46 & p_45_44;
 assign g_49_44 = g_49_46 | (p_49_46 & g_45_44);
 assign p_49_45 = p_49_46 & p_45_45;
 assign g_49_45 = g_49_46 | (p_49_46 & g_45_45);
 assign p_49_46 = p_49_48 & p_47_46;
 assign g_49_46 = g_49_48 | (p_49_48 & g_47_46);
 assign p_49_47 = p_49_48 & p_47_47;
 assign g_49_47 = g_49_48 | (p_49_48 & g_47_47);
 assign p_49_48 = p_49_49 & p_48_48;
 assign g_49_48 = g_49_49 | (p_49_49 & g_48_48);
 assign sum[49] = p_49_49^ g_48_0;
 assign p_50_0 = p_50_19 & p_18_0;
 assign g_50_0 = g_50_19 | (p_50_19 & g_18_0);
 assign p_50_1 = p_50_19 & p_18_1;
 assign g_50_1 = g_50_19 | (p_50_19 & g_18_1);
 assign p_50_2 = p_50_19 & p_18_2;
 assign g_50_2 = g_50_19 | (p_50_19 & g_18_2);
 assign p_50_3 = p_50_19 & p_18_3;
 assign g_50_3 = g_50_19 | (p_50_19 & g_18_3);
 assign p_50_4 = p_50_19 & p_18_4;
 assign g_50_4 = g_50_19 | (p_50_19 & g_18_4);
 assign p_50_5 = p_50_19 & p_18_5;
 assign g_50_5 = g_50_19 | (p_50_19 & g_18_5);
 assign p_50_6 = p_50_19 & p_18_6;
 assign g_50_6 = g_50_19 | (p_50_19 & g_18_6);
 assign p_50_7 = p_50_19 & p_18_7;
 assign g_50_7 = g_50_19 | (p_50_19 & g_18_7);
 assign p_50_8 = p_50_19 & p_18_8;
 assign g_50_8 = g_50_19 | (p_50_19 & g_18_8);
 assign p_50_9 = p_50_19 & p_18_9;
 assign g_50_9 = g_50_19 | (p_50_19 & g_18_9);
 assign p_50_10 = p_50_19 & p_18_10;
 assign g_50_10 = g_50_19 | (p_50_19 & g_18_10);
 assign p_50_11 = p_50_19 & p_18_11;
 assign g_50_11 = g_50_19 | (p_50_19 & g_18_11);
 assign p_50_12 = p_50_19 & p_18_12;
 assign g_50_12 = g_50_19 | (p_50_19 & g_18_12);
 assign p_50_13 = p_50_19 & p_18_13;
 assign g_50_13 = g_50_19 | (p_50_19 & g_18_13);
 assign p_50_14 = p_50_19 & p_18_14;
 assign g_50_14 = g_50_19 | (p_50_19 & g_18_14);
 assign p_50_15 = p_50_19 & p_18_15;
 assign g_50_15 = g_50_19 | (p_50_19 & g_18_15);
 assign p_50_16 = p_50_19 & p_18_16;
 assign g_50_16 = g_50_19 | (p_50_19 & g_18_16);
 assign p_50_17 = p_50_19 & p_18_17;
 assign g_50_17 = g_50_19 | (p_50_19 & g_18_17);
 assign p_50_18 = p_50_19 & p_18_18;
 assign g_50_18 = g_50_19 | (p_50_19 & g_18_18);
 assign p_50_19 = p_50_35 & p_34_19;
 assign g_50_19 = g_50_35 | (p_50_35 & g_34_19);
 assign p_50_20 = p_50_35 & p_34_20;
 assign g_50_20 = g_50_35 | (p_50_35 & g_34_20);
 assign p_50_21 = p_50_35 & p_34_21;
 assign g_50_21 = g_50_35 | (p_50_35 & g_34_21);
 assign p_50_22 = p_50_35 & p_34_22;
 assign g_50_22 = g_50_35 | (p_50_35 & g_34_22);
 assign p_50_23 = p_50_35 & p_34_23;
 assign g_50_23 = g_50_35 | (p_50_35 & g_34_23);
 assign p_50_24 = p_50_35 & p_34_24;
 assign g_50_24 = g_50_35 | (p_50_35 & g_34_24);
 assign p_50_25 = p_50_35 & p_34_25;
 assign g_50_25 = g_50_35 | (p_50_35 & g_34_25);
 assign p_50_26 = p_50_35 & p_34_26;
 assign g_50_26 = g_50_35 | (p_50_35 & g_34_26);
 assign p_50_27 = p_50_35 & p_34_27;
 assign g_50_27 = g_50_35 | (p_50_35 & g_34_27);
 assign p_50_28 = p_50_35 & p_34_28;
 assign g_50_28 = g_50_35 | (p_50_35 & g_34_28);
 assign p_50_29 = p_50_35 & p_34_29;
 assign g_50_29 = g_50_35 | (p_50_35 & g_34_29);
 assign p_50_30 = p_50_35 & p_34_30;
 assign g_50_30 = g_50_35 | (p_50_35 & g_34_30);
 assign p_50_31 = p_50_35 & p_34_31;
 assign g_50_31 = g_50_35 | (p_50_35 & g_34_31);
 assign p_50_32 = p_50_35 & p_34_32;
 assign g_50_32 = g_50_35 | (p_50_35 & g_34_32);
 assign p_50_33 = p_50_35 & p_34_33;
 assign g_50_33 = g_50_35 | (p_50_35 & g_34_33);
 assign p_50_34 = p_50_35 & p_34_34;
 assign g_50_34 = g_50_35 | (p_50_35 & g_34_34);
 assign p_50_35 = p_50_43 & p_42_35;
 assign g_50_35 = g_50_43 | (p_50_43 & g_42_35);
 assign p_50_36 = p_50_43 & p_42_36;
 assign g_50_36 = g_50_43 | (p_50_43 & g_42_36);
 assign p_50_37 = p_50_43 & p_42_37;
 assign g_50_37 = g_50_43 | (p_50_43 & g_42_37);
 assign p_50_38 = p_50_43 & p_42_38;
 assign g_50_38 = g_50_43 | (p_50_43 & g_42_38);
 assign p_50_39 = p_50_43 & p_42_39;
 assign g_50_39 = g_50_43 | (p_50_43 & g_42_39);
 assign p_50_40 = p_50_43 & p_42_40;
 assign g_50_40 = g_50_43 | (p_50_43 & g_42_40);
 assign p_50_41 = p_50_43 & p_42_41;
 assign g_50_41 = g_50_43 | (p_50_43 & g_42_41);
 assign p_50_42 = p_50_43 & p_42_42;
 assign g_50_42 = g_50_43 | (p_50_43 & g_42_42);
 assign p_50_43 = p_50_47 & p_46_43;
 assign g_50_43 = g_50_47 | (p_50_47 & g_46_43);
 assign p_50_44 = p_50_47 & p_46_44;
 assign g_50_44 = g_50_47 | (p_50_47 & g_46_44);
 assign p_50_45 = p_50_47 & p_46_45;
 assign g_50_45 = g_50_47 | (p_50_47 & g_46_45);
 assign p_50_46 = p_50_47 & p_46_46;
 assign g_50_46 = g_50_47 | (p_50_47 & g_46_46);
 assign p_50_47 = p_50_49 & p_48_47;
 assign g_50_47 = g_50_49 | (p_50_49 & g_48_47);
 assign p_50_48 = p_50_49 & p_48_48;
 assign g_50_48 = g_50_49 | (p_50_49 & g_48_48);
 assign p_50_49 = p_50_50 & p_49_49;
 assign g_50_49 = g_50_50 | (p_50_50 & g_49_49);
 assign sum[50] = p_50_50^ g_49_0;
 assign p_51_0 = p_51_20 & p_19_0;
 assign g_51_0 = g_51_20 | (p_51_20 & g_19_0);
 assign p_51_1 = p_51_20 & p_19_1;
 assign g_51_1 = g_51_20 | (p_51_20 & g_19_1);
 assign p_51_2 = p_51_20 & p_19_2;
 assign g_51_2 = g_51_20 | (p_51_20 & g_19_2);
 assign p_51_3 = p_51_20 & p_19_3;
 assign g_51_3 = g_51_20 | (p_51_20 & g_19_3);
 assign p_51_4 = p_51_20 & p_19_4;
 assign g_51_4 = g_51_20 | (p_51_20 & g_19_4);
 assign p_51_5 = p_51_20 & p_19_5;
 assign g_51_5 = g_51_20 | (p_51_20 & g_19_5);
 assign p_51_6 = p_51_20 & p_19_6;
 assign g_51_6 = g_51_20 | (p_51_20 & g_19_6);
 assign p_51_7 = p_51_20 & p_19_7;
 assign g_51_7 = g_51_20 | (p_51_20 & g_19_7);
 assign p_51_8 = p_51_20 & p_19_8;
 assign g_51_8 = g_51_20 | (p_51_20 & g_19_8);
 assign p_51_9 = p_51_20 & p_19_9;
 assign g_51_9 = g_51_20 | (p_51_20 & g_19_9);
 assign p_51_10 = p_51_20 & p_19_10;
 assign g_51_10 = g_51_20 | (p_51_20 & g_19_10);
 assign p_51_11 = p_51_20 & p_19_11;
 assign g_51_11 = g_51_20 | (p_51_20 & g_19_11);
 assign p_51_12 = p_51_20 & p_19_12;
 assign g_51_12 = g_51_20 | (p_51_20 & g_19_12);
 assign p_51_13 = p_51_20 & p_19_13;
 assign g_51_13 = g_51_20 | (p_51_20 & g_19_13);
 assign p_51_14 = p_51_20 & p_19_14;
 assign g_51_14 = g_51_20 | (p_51_20 & g_19_14);
 assign p_51_15 = p_51_20 & p_19_15;
 assign g_51_15 = g_51_20 | (p_51_20 & g_19_15);
 assign p_51_16 = p_51_20 & p_19_16;
 assign g_51_16 = g_51_20 | (p_51_20 & g_19_16);
 assign p_51_17 = p_51_20 & p_19_17;
 assign g_51_17 = g_51_20 | (p_51_20 & g_19_17);
 assign p_51_18 = p_51_20 & p_19_18;
 assign g_51_18 = g_51_20 | (p_51_20 & g_19_18);
 assign p_51_19 = p_51_20 & p_19_19;
 assign g_51_19 = g_51_20 | (p_51_20 & g_19_19);
 assign p_51_20 = p_51_36 & p_35_20;
 assign g_51_20 = g_51_36 | (p_51_36 & g_35_20);
 assign p_51_21 = p_51_36 & p_35_21;
 assign g_51_21 = g_51_36 | (p_51_36 & g_35_21);
 assign p_51_22 = p_51_36 & p_35_22;
 assign g_51_22 = g_51_36 | (p_51_36 & g_35_22);
 assign p_51_23 = p_51_36 & p_35_23;
 assign g_51_23 = g_51_36 | (p_51_36 & g_35_23);
 assign p_51_24 = p_51_36 & p_35_24;
 assign g_51_24 = g_51_36 | (p_51_36 & g_35_24);
 assign p_51_25 = p_51_36 & p_35_25;
 assign g_51_25 = g_51_36 | (p_51_36 & g_35_25);
 assign p_51_26 = p_51_36 & p_35_26;
 assign g_51_26 = g_51_36 | (p_51_36 & g_35_26);
 assign p_51_27 = p_51_36 & p_35_27;
 assign g_51_27 = g_51_36 | (p_51_36 & g_35_27);
 assign p_51_28 = p_51_36 & p_35_28;
 assign g_51_28 = g_51_36 | (p_51_36 & g_35_28);
 assign p_51_29 = p_51_36 & p_35_29;
 assign g_51_29 = g_51_36 | (p_51_36 & g_35_29);
 assign p_51_30 = p_51_36 & p_35_30;
 assign g_51_30 = g_51_36 | (p_51_36 & g_35_30);
 assign p_51_31 = p_51_36 & p_35_31;
 assign g_51_31 = g_51_36 | (p_51_36 & g_35_31);
 assign p_51_32 = p_51_36 & p_35_32;
 assign g_51_32 = g_51_36 | (p_51_36 & g_35_32);
 assign p_51_33 = p_51_36 & p_35_33;
 assign g_51_33 = g_51_36 | (p_51_36 & g_35_33);
 assign p_51_34 = p_51_36 & p_35_34;
 assign g_51_34 = g_51_36 | (p_51_36 & g_35_34);
 assign p_51_35 = p_51_36 & p_35_35;
 assign g_51_35 = g_51_36 | (p_51_36 & g_35_35);
 assign p_51_36 = p_51_44 & p_43_36;
 assign g_51_36 = g_51_44 | (p_51_44 & g_43_36);
 assign p_51_37 = p_51_44 & p_43_37;
 assign g_51_37 = g_51_44 | (p_51_44 & g_43_37);
 assign p_51_38 = p_51_44 & p_43_38;
 assign g_51_38 = g_51_44 | (p_51_44 & g_43_38);
 assign p_51_39 = p_51_44 & p_43_39;
 assign g_51_39 = g_51_44 | (p_51_44 & g_43_39);
 assign p_51_40 = p_51_44 & p_43_40;
 assign g_51_40 = g_51_44 | (p_51_44 & g_43_40);
 assign p_51_41 = p_51_44 & p_43_41;
 assign g_51_41 = g_51_44 | (p_51_44 & g_43_41);
 assign p_51_42 = p_51_44 & p_43_42;
 assign g_51_42 = g_51_44 | (p_51_44 & g_43_42);
 assign p_51_43 = p_51_44 & p_43_43;
 assign g_51_43 = g_51_44 | (p_51_44 & g_43_43);
 assign p_51_44 = p_51_48 & p_47_44;
 assign g_51_44 = g_51_48 | (p_51_48 & g_47_44);
 assign p_51_45 = p_51_48 & p_47_45;
 assign g_51_45 = g_51_48 | (p_51_48 & g_47_45);
 assign p_51_46 = p_51_48 & p_47_46;
 assign g_51_46 = g_51_48 | (p_51_48 & g_47_46);
 assign p_51_47 = p_51_48 & p_47_47;
 assign g_51_47 = g_51_48 | (p_51_48 & g_47_47);
 assign p_51_48 = p_51_50 & p_49_48;
 assign g_51_48 = g_51_50 | (p_51_50 & g_49_48);
 assign p_51_49 = p_51_50 & p_49_49;
 assign g_51_49 = g_51_50 | (p_51_50 & g_49_49);
 assign p_51_50 = p_51_51 & p_50_50;
 assign g_51_50 = g_51_51 | (p_51_51 & g_50_50);
 assign sum[51] = p_51_51^ g_50_0;
 assign p_52_0 = p_52_21 & p_20_0;
 assign g_52_0 = g_52_21 | (p_52_21 & g_20_0);
 assign p_52_1 = p_52_21 & p_20_1;
 assign g_52_1 = g_52_21 | (p_52_21 & g_20_1);
 assign p_52_2 = p_52_21 & p_20_2;
 assign g_52_2 = g_52_21 | (p_52_21 & g_20_2);
 assign p_52_3 = p_52_21 & p_20_3;
 assign g_52_3 = g_52_21 | (p_52_21 & g_20_3);
 assign p_52_4 = p_52_21 & p_20_4;
 assign g_52_4 = g_52_21 | (p_52_21 & g_20_4);
 assign p_52_5 = p_52_21 & p_20_5;
 assign g_52_5 = g_52_21 | (p_52_21 & g_20_5);
 assign p_52_6 = p_52_21 & p_20_6;
 assign g_52_6 = g_52_21 | (p_52_21 & g_20_6);
 assign p_52_7 = p_52_21 & p_20_7;
 assign g_52_7 = g_52_21 | (p_52_21 & g_20_7);
 assign p_52_8 = p_52_21 & p_20_8;
 assign g_52_8 = g_52_21 | (p_52_21 & g_20_8);
 assign p_52_9 = p_52_21 & p_20_9;
 assign g_52_9 = g_52_21 | (p_52_21 & g_20_9);
 assign p_52_10 = p_52_21 & p_20_10;
 assign g_52_10 = g_52_21 | (p_52_21 & g_20_10);
 assign p_52_11 = p_52_21 & p_20_11;
 assign g_52_11 = g_52_21 | (p_52_21 & g_20_11);
 assign p_52_12 = p_52_21 & p_20_12;
 assign g_52_12 = g_52_21 | (p_52_21 & g_20_12);
 assign p_52_13 = p_52_21 & p_20_13;
 assign g_52_13 = g_52_21 | (p_52_21 & g_20_13);
 assign p_52_14 = p_52_21 & p_20_14;
 assign g_52_14 = g_52_21 | (p_52_21 & g_20_14);
 assign p_52_15 = p_52_21 & p_20_15;
 assign g_52_15 = g_52_21 | (p_52_21 & g_20_15);
 assign p_52_16 = p_52_21 & p_20_16;
 assign g_52_16 = g_52_21 | (p_52_21 & g_20_16);
 assign p_52_17 = p_52_21 & p_20_17;
 assign g_52_17 = g_52_21 | (p_52_21 & g_20_17);
 assign p_52_18 = p_52_21 & p_20_18;
 assign g_52_18 = g_52_21 | (p_52_21 & g_20_18);
 assign p_52_19 = p_52_21 & p_20_19;
 assign g_52_19 = g_52_21 | (p_52_21 & g_20_19);
 assign p_52_20 = p_52_21 & p_20_20;
 assign g_52_20 = g_52_21 | (p_52_21 & g_20_20);
 assign p_52_21 = p_52_37 & p_36_21;
 assign g_52_21 = g_52_37 | (p_52_37 & g_36_21);
 assign p_52_22 = p_52_37 & p_36_22;
 assign g_52_22 = g_52_37 | (p_52_37 & g_36_22);
 assign p_52_23 = p_52_37 & p_36_23;
 assign g_52_23 = g_52_37 | (p_52_37 & g_36_23);
 assign p_52_24 = p_52_37 & p_36_24;
 assign g_52_24 = g_52_37 | (p_52_37 & g_36_24);
 assign p_52_25 = p_52_37 & p_36_25;
 assign g_52_25 = g_52_37 | (p_52_37 & g_36_25);
 assign p_52_26 = p_52_37 & p_36_26;
 assign g_52_26 = g_52_37 | (p_52_37 & g_36_26);
 assign p_52_27 = p_52_37 & p_36_27;
 assign g_52_27 = g_52_37 | (p_52_37 & g_36_27);
 assign p_52_28 = p_52_37 & p_36_28;
 assign g_52_28 = g_52_37 | (p_52_37 & g_36_28);
 assign p_52_29 = p_52_37 & p_36_29;
 assign g_52_29 = g_52_37 | (p_52_37 & g_36_29);
 assign p_52_30 = p_52_37 & p_36_30;
 assign g_52_30 = g_52_37 | (p_52_37 & g_36_30);
 assign p_52_31 = p_52_37 & p_36_31;
 assign g_52_31 = g_52_37 | (p_52_37 & g_36_31);
 assign p_52_32 = p_52_37 & p_36_32;
 assign g_52_32 = g_52_37 | (p_52_37 & g_36_32);
 assign p_52_33 = p_52_37 & p_36_33;
 assign g_52_33 = g_52_37 | (p_52_37 & g_36_33);
 assign p_52_34 = p_52_37 & p_36_34;
 assign g_52_34 = g_52_37 | (p_52_37 & g_36_34);
 assign p_52_35 = p_52_37 & p_36_35;
 assign g_52_35 = g_52_37 | (p_52_37 & g_36_35);
 assign p_52_36 = p_52_37 & p_36_36;
 assign g_52_36 = g_52_37 | (p_52_37 & g_36_36);
 assign p_52_37 = p_52_45 & p_44_37;
 assign g_52_37 = g_52_45 | (p_52_45 & g_44_37);
 assign p_52_38 = p_52_45 & p_44_38;
 assign g_52_38 = g_52_45 | (p_52_45 & g_44_38);
 assign p_52_39 = p_52_45 & p_44_39;
 assign g_52_39 = g_52_45 | (p_52_45 & g_44_39);
 assign p_52_40 = p_52_45 & p_44_40;
 assign g_52_40 = g_52_45 | (p_52_45 & g_44_40);
 assign p_52_41 = p_52_45 & p_44_41;
 assign g_52_41 = g_52_45 | (p_52_45 & g_44_41);
 assign p_52_42 = p_52_45 & p_44_42;
 assign g_52_42 = g_52_45 | (p_52_45 & g_44_42);
 assign p_52_43 = p_52_45 & p_44_43;
 assign g_52_43 = g_52_45 | (p_52_45 & g_44_43);
 assign p_52_44 = p_52_45 & p_44_44;
 assign g_52_44 = g_52_45 | (p_52_45 & g_44_44);
 assign p_52_45 = p_52_49 & p_48_45;
 assign g_52_45 = g_52_49 | (p_52_49 & g_48_45);
 assign p_52_46 = p_52_49 & p_48_46;
 assign g_52_46 = g_52_49 | (p_52_49 & g_48_46);
 assign p_52_47 = p_52_49 & p_48_47;
 assign g_52_47 = g_52_49 | (p_52_49 & g_48_47);
 assign p_52_48 = p_52_49 & p_48_48;
 assign g_52_48 = g_52_49 | (p_52_49 & g_48_48);
 assign p_52_49 = p_52_51 & p_50_49;
 assign g_52_49 = g_52_51 | (p_52_51 & g_50_49);
 assign p_52_50 = p_52_51 & p_50_50;
 assign g_52_50 = g_52_51 | (p_52_51 & g_50_50);
 assign p_52_51 = p_52_52 & p_51_51;
 assign g_52_51 = g_52_52 | (p_52_52 & g_51_51);
 assign sum[52] = p_52_52^ g_51_0;
 assign p_53_0 = p_53_22 & p_21_0;
 assign g_53_0 = g_53_22 | (p_53_22 & g_21_0);
 assign p_53_1 = p_53_22 & p_21_1;
 assign g_53_1 = g_53_22 | (p_53_22 & g_21_1);
 assign p_53_2 = p_53_22 & p_21_2;
 assign g_53_2 = g_53_22 | (p_53_22 & g_21_2);
 assign p_53_3 = p_53_22 & p_21_3;
 assign g_53_3 = g_53_22 | (p_53_22 & g_21_3);
 assign p_53_4 = p_53_22 & p_21_4;
 assign g_53_4 = g_53_22 | (p_53_22 & g_21_4);
 assign p_53_5 = p_53_22 & p_21_5;
 assign g_53_5 = g_53_22 | (p_53_22 & g_21_5);
 assign p_53_6 = p_53_22 & p_21_6;
 assign g_53_6 = g_53_22 | (p_53_22 & g_21_6);
 assign p_53_7 = p_53_22 & p_21_7;
 assign g_53_7 = g_53_22 | (p_53_22 & g_21_7);
 assign p_53_8 = p_53_22 & p_21_8;
 assign g_53_8 = g_53_22 | (p_53_22 & g_21_8);
 assign p_53_9 = p_53_22 & p_21_9;
 assign g_53_9 = g_53_22 | (p_53_22 & g_21_9);
 assign p_53_10 = p_53_22 & p_21_10;
 assign g_53_10 = g_53_22 | (p_53_22 & g_21_10);
 assign p_53_11 = p_53_22 & p_21_11;
 assign g_53_11 = g_53_22 | (p_53_22 & g_21_11);
 assign p_53_12 = p_53_22 & p_21_12;
 assign g_53_12 = g_53_22 | (p_53_22 & g_21_12);
 assign p_53_13 = p_53_22 & p_21_13;
 assign g_53_13 = g_53_22 | (p_53_22 & g_21_13);
 assign p_53_14 = p_53_22 & p_21_14;
 assign g_53_14 = g_53_22 | (p_53_22 & g_21_14);
 assign p_53_15 = p_53_22 & p_21_15;
 assign g_53_15 = g_53_22 | (p_53_22 & g_21_15);
 assign p_53_16 = p_53_22 & p_21_16;
 assign g_53_16 = g_53_22 | (p_53_22 & g_21_16);
 assign p_53_17 = p_53_22 & p_21_17;
 assign g_53_17 = g_53_22 | (p_53_22 & g_21_17);
 assign p_53_18 = p_53_22 & p_21_18;
 assign g_53_18 = g_53_22 | (p_53_22 & g_21_18);
 assign p_53_19 = p_53_22 & p_21_19;
 assign g_53_19 = g_53_22 | (p_53_22 & g_21_19);
 assign p_53_20 = p_53_22 & p_21_20;
 assign g_53_20 = g_53_22 | (p_53_22 & g_21_20);
 assign p_53_21 = p_53_22 & p_21_21;
 assign g_53_21 = g_53_22 | (p_53_22 & g_21_21);
 assign p_53_22 = p_53_38 & p_37_22;
 assign g_53_22 = g_53_38 | (p_53_38 & g_37_22);
 assign p_53_23 = p_53_38 & p_37_23;
 assign g_53_23 = g_53_38 | (p_53_38 & g_37_23);
 assign p_53_24 = p_53_38 & p_37_24;
 assign g_53_24 = g_53_38 | (p_53_38 & g_37_24);
 assign p_53_25 = p_53_38 & p_37_25;
 assign g_53_25 = g_53_38 | (p_53_38 & g_37_25);
 assign p_53_26 = p_53_38 & p_37_26;
 assign g_53_26 = g_53_38 | (p_53_38 & g_37_26);
 assign p_53_27 = p_53_38 & p_37_27;
 assign g_53_27 = g_53_38 | (p_53_38 & g_37_27);
 assign p_53_28 = p_53_38 & p_37_28;
 assign g_53_28 = g_53_38 | (p_53_38 & g_37_28);
 assign p_53_29 = p_53_38 & p_37_29;
 assign g_53_29 = g_53_38 | (p_53_38 & g_37_29);
 assign p_53_30 = p_53_38 & p_37_30;
 assign g_53_30 = g_53_38 | (p_53_38 & g_37_30);
 assign p_53_31 = p_53_38 & p_37_31;
 assign g_53_31 = g_53_38 | (p_53_38 & g_37_31);
 assign p_53_32 = p_53_38 & p_37_32;
 assign g_53_32 = g_53_38 | (p_53_38 & g_37_32);
 assign p_53_33 = p_53_38 & p_37_33;
 assign g_53_33 = g_53_38 | (p_53_38 & g_37_33);
 assign p_53_34 = p_53_38 & p_37_34;
 assign g_53_34 = g_53_38 | (p_53_38 & g_37_34);
 assign p_53_35 = p_53_38 & p_37_35;
 assign g_53_35 = g_53_38 | (p_53_38 & g_37_35);
 assign p_53_36 = p_53_38 & p_37_36;
 assign g_53_36 = g_53_38 | (p_53_38 & g_37_36);
 assign p_53_37 = p_53_38 & p_37_37;
 assign g_53_37 = g_53_38 | (p_53_38 & g_37_37);
 assign p_53_38 = p_53_46 & p_45_38;
 assign g_53_38 = g_53_46 | (p_53_46 & g_45_38);
 assign p_53_39 = p_53_46 & p_45_39;
 assign g_53_39 = g_53_46 | (p_53_46 & g_45_39);
 assign p_53_40 = p_53_46 & p_45_40;
 assign g_53_40 = g_53_46 | (p_53_46 & g_45_40);
 assign p_53_41 = p_53_46 & p_45_41;
 assign g_53_41 = g_53_46 | (p_53_46 & g_45_41);
 assign p_53_42 = p_53_46 & p_45_42;
 assign g_53_42 = g_53_46 | (p_53_46 & g_45_42);
 assign p_53_43 = p_53_46 & p_45_43;
 assign g_53_43 = g_53_46 | (p_53_46 & g_45_43);
 assign p_53_44 = p_53_46 & p_45_44;
 assign g_53_44 = g_53_46 | (p_53_46 & g_45_44);
 assign p_53_45 = p_53_46 & p_45_45;
 assign g_53_45 = g_53_46 | (p_53_46 & g_45_45);
 assign p_53_46 = p_53_50 & p_49_46;
 assign g_53_46 = g_53_50 | (p_53_50 & g_49_46);
 assign p_53_47 = p_53_50 & p_49_47;
 assign g_53_47 = g_53_50 | (p_53_50 & g_49_47);
 assign p_53_48 = p_53_50 & p_49_48;
 assign g_53_48 = g_53_50 | (p_53_50 & g_49_48);
 assign p_53_49 = p_53_50 & p_49_49;
 assign g_53_49 = g_53_50 | (p_53_50 & g_49_49);
 assign p_53_50 = p_53_52 & p_51_50;
 assign g_53_50 = g_53_52 | (p_53_52 & g_51_50);
 assign p_53_51 = p_53_52 & p_51_51;
 assign g_53_51 = g_53_52 | (p_53_52 & g_51_51);
 assign p_53_52 = p_53_53 & p_52_52;
 assign g_53_52 = g_53_53 | (p_53_53 & g_52_52);
 assign sum[53] = p_53_53^ g_52_0;
 assign p_54_0 = p_54_23 & p_22_0;
 assign g_54_0 = g_54_23 | (p_54_23 & g_22_0);
 assign p_54_1 = p_54_23 & p_22_1;
 assign g_54_1 = g_54_23 | (p_54_23 & g_22_1);
 assign p_54_2 = p_54_23 & p_22_2;
 assign g_54_2 = g_54_23 | (p_54_23 & g_22_2);
 assign p_54_3 = p_54_23 & p_22_3;
 assign g_54_3 = g_54_23 | (p_54_23 & g_22_3);
 assign p_54_4 = p_54_23 & p_22_4;
 assign g_54_4 = g_54_23 | (p_54_23 & g_22_4);
 assign p_54_5 = p_54_23 & p_22_5;
 assign g_54_5 = g_54_23 | (p_54_23 & g_22_5);
 assign p_54_6 = p_54_23 & p_22_6;
 assign g_54_6 = g_54_23 | (p_54_23 & g_22_6);
 assign p_54_7 = p_54_23 & p_22_7;
 assign g_54_7 = g_54_23 | (p_54_23 & g_22_7);
 assign p_54_8 = p_54_23 & p_22_8;
 assign g_54_8 = g_54_23 | (p_54_23 & g_22_8);
 assign p_54_9 = p_54_23 & p_22_9;
 assign g_54_9 = g_54_23 | (p_54_23 & g_22_9);
 assign p_54_10 = p_54_23 & p_22_10;
 assign g_54_10 = g_54_23 | (p_54_23 & g_22_10);
 assign p_54_11 = p_54_23 & p_22_11;
 assign g_54_11 = g_54_23 | (p_54_23 & g_22_11);
 assign p_54_12 = p_54_23 & p_22_12;
 assign g_54_12 = g_54_23 | (p_54_23 & g_22_12);
 assign p_54_13 = p_54_23 & p_22_13;
 assign g_54_13 = g_54_23 | (p_54_23 & g_22_13);
 assign p_54_14 = p_54_23 & p_22_14;
 assign g_54_14 = g_54_23 | (p_54_23 & g_22_14);
 assign p_54_15 = p_54_23 & p_22_15;
 assign g_54_15 = g_54_23 | (p_54_23 & g_22_15);
 assign p_54_16 = p_54_23 & p_22_16;
 assign g_54_16 = g_54_23 | (p_54_23 & g_22_16);
 assign p_54_17 = p_54_23 & p_22_17;
 assign g_54_17 = g_54_23 | (p_54_23 & g_22_17);
 assign p_54_18 = p_54_23 & p_22_18;
 assign g_54_18 = g_54_23 | (p_54_23 & g_22_18);
 assign p_54_19 = p_54_23 & p_22_19;
 assign g_54_19 = g_54_23 | (p_54_23 & g_22_19);
 assign p_54_20 = p_54_23 & p_22_20;
 assign g_54_20 = g_54_23 | (p_54_23 & g_22_20);
 assign p_54_21 = p_54_23 & p_22_21;
 assign g_54_21 = g_54_23 | (p_54_23 & g_22_21);
 assign p_54_22 = p_54_23 & p_22_22;
 assign g_54_22 = g_54_23 | (p_54_23 & g_22_22);
 assign p_54_23 = p_54_39 & p_38_23;
 assign g_54_23 = g_54_39 | (p_54_39 & g_38_23);
 assign p_54_24 = p_54_39 & p_38_24;
 assign g_54_24 = g_54_39 | (p_54_39 & g_38_24);
 assign p_54_25 = p_54_39 & p_38_25;
 assign g_54_25 = g_54_39 | (p_54_39 & g_38_25);
 assign p_54_26 = p_54_39 & p_38_26;
 assign g_54_26 = g_54_39 | (p_54_39 & g_38_26);
 assign p_54_27 = p_54_39 & p_38_27;
 assign g_54_27 = g_54_39 | (p_54_39 & g_38_27);
 assign p_54_28 = p_54_39 & p_38_28;
 assign g_54_28 = g_54_39 | (p_54_39 & g_38_28);
 assign p_54_29 = p_54_39 & p_38_29;
 assign g_54_29 = g_54_39 | (p_54_39 & g_38_29);
 assign p_54_30 = p_54_39 & p_38_30;
 assign g_54_30 = g_54_39 | (p_54_39 & g_38_30);
 assign p_54_31 = p_54_39 & p_38_31;
 assign g_54_31 = g_54_39 | (p_54_39 & g_38_31);
 assign p_54_32 = p_54_39 & p_38_32;
 assign g_54_32 = g_54_39 | (p_54_39 & g_38_32);
 assign p_54_33 = p_54_39 & p_38_33;
 assign g_54_33 = g_54_39 | (p_54_39 & g_38_33);
 assign p_54_34 = p_54_39 & p_38_34;
 assign g_54_34 = g_54_39 | (p_54_39 & g_38_34);
 assign p_54_35 = p_54_39 & p_38_35;
 assign g_54_35 = g_54_39 | (p_54_39 & g_38_35);
 assign p_54_36 = p_54_39 & p_38_36;
 assign g_54_36 = g_54_39 | (p_54_39 & g_38_36);
 assign p_54_37 = p_54_39 & p_38_37;
 assign g_54_37 = g_54_39 | (p_54_39 & g_38_37);
 assign p_54_38 = p_54_39 & p_38_38;
 assign g_54_38 = g_54_39 | (p_54_39 & g_38_38);
 assign p_54_39 = p_54_47 & p_46_39;
 assign g_54_39 = g_54_47 | (p_54_47 & g_46_39);
 assign p_54_40 = p_54_47 & p_46_40;
 assign g_54_40 = g_54_47 | (p_54_47 & g_46_40);
 assign p_54_41 = p_54_47 & p_46_41;
 assign g_54_41 = g_54_47 | (p_54_47 & g_46_41);
 assign p_54_42 = p_54_47 & p_46_42;
 assign g_54_42 = g_54_47 | (p_54_47 & g_46_42);
 assign p_54_43 = p_54_47 & p_46_43;
 assign g_54_43 = g_54_47 | (p_54_47 & g_46_43);
 assign p_54_44 = p_54_47 & p_46_44;
 assign g_54_44 = g_54_47 | (p_54_47 & g_46_44);
 assign p_54_45 = p_54_47 & p_46_45;
 assign g_54_45 = g_54_47 | (p_54_47 & g_46_45);
 assign p_54_46 = p_54_47 & p_46_46;
 assign g_54_46 = g_54_47 | (p_54_47 & g_46_46);
 assign p_54_47 = p_54_51 & p_50_47;
 assign g_54_47 = g_54_51 | (p_54_51 & g_50_47);
 assign p_54_48 = p_54_51 & p_50_48;
 assign g_54_48 = g_54_51 | (p_54_51 & g_50_48);
 assign p_54_49 = p_54_51 & p_50_49;
 assign g_54_49 = g_54_51 | (p_54_51 & g_50_49);
 assign p_54_50 = p_54_51 & p_50_50;
 assign g_54_50 = g_54_51 | (p_54_51 & g_50_50);
 assign p_54_51 = p_54_53 & p_52_51;
 assign g_54_51 = g_54_53 | (p_54_53 & g_52_51);
 assign p_54_52 = p_54_53 & p_52_52;
 assign g_54_52 = g_54_53 | (p_54_53 & g_52_52);
 assign p_54_53 = p_54_54 & p_53_53;
 assign g_54_53 = g_54_54 | (p_54_54 & g_53_53);
 assign sum[54] = p_54_54^ g_53_0;
 assign p_55_0 = p_55_24 & p_23_0;
 assign g_55_0 = g_55_24 | (p_55_24 & g_23_0);
 assign p_55_1 = p_55_24 & p_23_1;
 assign g_55_1 = g_55_24 | (p_55_24 & g_23_1);
 assign p_55_2 = p_55_24 & p_23_2;
 assign g_55_2 = g_55_24 | (p_55_24 & g_23_2);
 assign p_55_3 = p_55_24 & p_23_3;
 assign g_55_3 = g_55_24 | (p_55_24 & g_23_3);
 assign p_55_4 = p_55_24 & p_23_4;
 assign g_55_4 = g_55_24 | (p_55_24 & g_23_4);
 assign p_55_5 = p_55_24 & p_23_5;
 assign g_55_5 = g_55_24 | (p_55_24 & g_23_5);
 assign p_55_6 = p_55_24 & p_23_6;
 assign g_55_6 = g_55_24 | (p_55_24 & g_23_6);
 assign p_55_7 = p_55_24 & p_23_7;
 assign g_55_7 = g_55_24 | (p_55_24 & g_23_7);
 assign p_55_8 = p_55_24 & p_23_8;
 assign g_55_8 = g_55_24 | (p_55_24 & g_23_8);
 assign p_55_9 = p_55_24 & p_23_9;
 assign g_55_9 = g_55_24 | (p_55_24 & g_23_9);
 assign p_55_10 = p_55_24 & p_23_10;
 assign g_55_10 = g_55_24 | (p_55_24 & g_23_10);
 assign p_55_11 = p_55_24 & p_23_11;
 assign g_55_11 = g_55_24 | (p_55_24 & g_23_11);
 assign p_55_12 = p_55_24 & p_23_12;
 assign g_55_12 = g_55_24 | (p_55_24 & g_23_12);
 assign p_55_13 = p_55_24 & p_23_13;
 assign g_55_13 = g_55_24 | (p_55_24 & g_23_13);
 assign p_55_14 = p_55_24 & p_23_14;
 assign g_55_14 = g_55_24 | (p_55_24 & g_23_14);
 assign p_55_15 = p_55_24 & p_23_15;
 assign g_55_15 = g_55_24 | (p_55_24 & g_23_15);
 assign p_55_16 = p_55_24 & p_23_16;
 assign g_55_16 = g_55_24 | (p_55_24 & g_23_16);
 assign p_55_17 = p_55_24 & p_23_17;
 assign g_55_17 = g_55_24 | (p_55_24 & g_23_17);
 assign p_55_18 = p_55_24 & p_23_18;
 assign g_55_18 = g_55_24 | (p_55_24 & g_23_18);
 assign p_55_19 = p_55_24 & p_23_19;
 assign g_55_19 = g_55_24 | (p_55_24 & g_23_19);
 assign p_55_20 = p_55_24 & p_23_20;
 assign g_55_20 = g_55_24 | (p_55_24 & g_23_20);
 assign p_55_21 = p_55_24 & p_23_21;
 assign g_55_21 = g_55_24 | (p_55_24 & g_23_21);
 assign p_55_22 = p_55_24 & p_23_22;
 assign g_55_22 = g_55_24 | (p_55_24 & g_23_22);
 assign p_55_23 = p_55_24 & p_23_23;
 assign g_55_23 = g_55_24 | (p_55_24 & g_23_23);
 assign p_55_24 = p_55_40 & p_39_24;
 assign g_55_24 = g_55_40 | (p_55_40 & g_39_24);
 assign p_55_25 = p_55_40 & p_39_25;
 assign g_55_25 = g_55_40 | (p_55_40 & g_39_25);
 assign p_55_26 = p_55_40 & p_39_26;
 assign g_55_26 = g_55_40 | (p_55_40 & g_39_26);
 assign p_55_27 = p_55_40 & p_39_27;
 assign g_55_27 = g_55_40 | (p_55_40 & g_39_27);
 assign p_55_28 = p_55_40 & p_39_28;
 assign g_55_28 = g_55_40 | (p_55_40 & g_39_28);
 assign p_55_29 = p_55_40 & p_39_29;
 assign g_55_29 = g_55_40 | (p_55_40 & g_39_29);
 assign p_55_30 = p_55_40 & p_39_30;
 assign g_55_30 = g_55_40 | (p_55_40 & g_39_30);
 assign p_55_31 = p_55_40 & p_39_31;
 assign g_55_31 = g_55_40 | (p_55_40 & g_39_31);
 assign p_55_32 = p_55_40 & p_39_32;
 assign g_55_32 = g_55_40 | (p_55_40 & g_39_32);
 assign p_55_33 = p_55_40 & p_39_33;
 assign g_55_33 = g_55_40 | (p_55_40 & g_39_33);
 assign p_55_34 = p_55_40 & p_39_34;
 assign g_55_34 = g_55_40 | (p_55_40 & g_39_34);
 assign p_55_35 = p_55_40 & p_39_35;
 assign g_55_35 = g_55_40 | (p_55_40 & g_39_35);
 assign p_55_36 = p_55_40 & p_39_36;
 assign g_55_36 = g_55_40 | (p_55_40 & g_39_36);
 assign p_55_37 = p_55_40 & p_39_37;
 assign g_55_37 = g_55_40 | (p_55_40 & g_39_37);
 assign p_55_38 = p_55_40 & p_39_38;
 assign g_55_38 = g_55_40 | (p_55_40 & g_39_38);
 assign p_55_39 = p_55_40 & p_39_39;
 assign g_55_39 = g_55_40 | (p_55_40 & g_39_39);
 assign p_55_40 = p_55_48 & p_47_40;
 assign g_55_40 = g_55_48 | (p_55_48 & g_47_40);
 assign p_55_41 = p_55_48 & p_47_41;
 assign g_55_41 = g_55_48 | (p_55_48 & g_47_41);
 assign p_55_42 = p_55_48 & p_47_42;
 assign g_55_42 = g_55_48 | (p_55_48 & g_47_42);
 assign p_55_43 = p_55_48 & p_47_43;
 assign g_55_43 = g_55_48 | (p_55_48 & g_47_43);
 assign p_55_44 = p_55_48 & p_47_44;
 assign g_55_44 = g_55_48 | (p_55_48 & g_47_44);
 assign p_55_45 = p_55_48 & p_47_45;
 assign g_55_45 = g_55_48 | (p_55_48 & g_47_45);
 assign p_55_46 = p_55_48 & p_47_46;
 assign g_55_46 = g_55_48 | (p_55_48 & g_47_46);
 assign p_55_47 = p_55_48 & p_47_47;
 assign g_55_47 = g_55_48 | (p_55_48 & g_47_47);
 assign p_55_48 = p_55_52 & p_51_48;
 assign g_55_48 = g_55_52 | (p_55_52 & g_51_48);
 assign p_55_49 = p_55_52 & p_51_49;
 assign g_55_49 = g_55_52 | (p_55_52 & g_51_49);
 assign p_55_50 = p_55_52 & p_51_50;
 assign g_55_50 = g_55_52 | (p_55_52 & g_51_50);
 assign p_55_51 = p_55_52 & p_51_51;
 assign g_55_51 = g_55_52 | (p_55_52 & g_51_51);
 assign p_55_52 = p_55_54 & p_53_52;
 assign g_55_52 = g_55_54 | (p_55_54 & g_53_52);
 assign p_55_53 = p_55_54 & p_53_53;
 assign g_55_53 = g_55_54 | (p_55_54 & g_53_53);
 assign p_55_54 = p_55_55 & p_54_54;
 assign g_55_54 = g_55_55 | (p_55_55 & g_54_54);
 assign sum[55] = p_55_55^ g_54_0;
 assign p_56_0 = p_56_25 & p_24_0;
 assign g_56_0 = g_56_25 | (p_56_25 & g_24_0);
 assign p_56_1 = p_56_25 & p_24_1;
 assign g_56_1 = g_56_25 | (p_56_25 & g_24_1);
 assign p_56_2 = p_56_25 & p_24_2;
 assign g_56_2 = g_56_25 | (p_56_25 & g_24_2);
 assign p_56_3 = p_56_25 & p_24_3;
 assign g_56_3 = g_56_25 | (p_56_25 & g_24_3);
 assign p_56_4 = p_56_25 & p_24_4;
 assign g_56_4 = g_56_25 | (p_56_25 & g_24_4);
 assign p_56_5 = p_56_25 & p_24_5;
 assign g_56_5 = g_56_25 | (p_56_25 & g_24_5);
 assign p_56_6 = p_56_25 & p_24_6;
 assign g_56_6 = g_56_25 | (p_56_25 & g_24_6);
 assign p_56_7 = p_56_25 & p_24_7;
 assign g_56_7 = g_56_25 | (p_56_25 & g_24_7);
 assign p_56_8 = p_56_25 & p_24_8;
 assign g_56_8 = g_56_25 | (p_56_25 & g_24_8);
 assign p_56_9 = p_56_25 & p_24_9;
 assign g_56_9 = g_56_25 | (p_56_25 & g_24_9);
 assign p_56_10 = p_56_25 & p_24_10;
 assign g_56_10 = g_56_25 | (p_56_25 & g_24_10);
 assign p_56_11 = p_56_25 & p_24_11;
 assign g_56_11 = g_56_25 | (p_56_25 & g_24_11);
 assign p_56_12 = p_56_25 & p_24_12;
 assign g_56_12 = g_56_25 | (p_56_25 & g_24_12);
 assign p_56_13 = p_56_25 & p_24_13;
 assign g_56_13 = g_56_25 | (p_56_25 & g_24_13);
 assign p_56_14 = p_56_25 & p_24_14;
 assign g_56_14 = g_56_25 | (p_56_25 & g_24_14);
 assign p_56_15 = p_56_25 & p_24_15;
 assign g_56_15 = g_56_25 | (p_56_25 & g_24_15);
 assign p_56_16 = p_56_25 & p_24_16;
 assign g_56_16 = g_56_25 | (p_56_25 & g_24_16);
 assign p_56_17 = p_56_25 & p_24_17;
 assign g_56_17 = g_56_25 | (p_56_25 & g_24_17);
 assign p_56_18 = p_56_25 & p_24_18;
 assign g_56_18 = g_56_25 | (p_56_25 & g_24_18);
 assign p_56_19 = p_56_25 & p_24_19;
 assign g_56_19 = g_56_25 | (p_56_25 & g_24_19);
 assign p_56_20 = p_56_25 & p_24_20;
 assign g_56_20 = g_56_25 | (p_56_25 & g_24_20);
 assign p_56_21 = p_56_25 & p_24_21;
 assign g_56_21 = g_56_25 | (p_56_25 & g_24_21);
 assign p_56_22 = p_56_25 & p_24_22;
 assign g_56_22 = g_56_25 | (p_56_25 & g_24_22);
 assign p_56_23 = p_56_25 & p_24_23;
 assign g_56_23 = g_56_25 | (p_56_25 & g_24_23);
 assign p_56_24 = p_56_25 & p_24_24;
 assign g_56_24 = g_56_25 | (p_56_25 & g_24_24);
 assign p_56_25 = p_56_41 & p_40_25;
 assign g_56_25 = g_56_41 | (p_56_41 & g_40_25);
 assign p_56_26 = p_56_41 & p_40_26;
 assign g_56_26 = g_56_41 | (p_56_41 & g_40_26);
 assign p_56_27 = p_56_41 & p_40_27;
 assign g_56_27 = g_56_41 | (p_56_41 & g_40_27);
 assign p_56_28 = p_56_41 & p_40_28;
 assign g_56_28 = g_56_41 | (p_56_41 & g_40_28);
 assign p_56_29 = p_56_41 & p_40_29;
 assign g_56_29 = g_56_41 | (p_56_41 & g_40_29);
 assign p_56_30 = p_56_41 & p_40_30;
 assign g_56_30 = g_56_41 | (p_56_41 & g_40_30);
 assign p_56_31 = p_56_41 & p_40_31;
 assign g_56_31 = g_56_41 | (p_56_41 & g_40_31);
 assign p_56_32 = p_56_41 & p_40_32;
 assign g_56_32 = g_56_41 | (p_56_41 & g_40_32);
 assign p_56_33 = p_56_41 & p_40_33;
 assign g_56_33 = g_56_41 | (p_56_41 & g_40_33);
 assign p_56_34 = p_56_41 & p_40_34;
 assign g_56_34 = g_56_41 | (p_56_41 & g_40_34);
 assign p_56_35 = p_56_41 & p_40_35;
 assign g_56_35 = g_56_41 | (p_56_41 & g_40_35);
 assign p_56_36 = p_56_41 & p_40_36;
 assign g_56_36 = g_56_41 | (p_56_41 & g_40_36);
 assign p_56_37 = p_56_41 & p_40_37;
 assign g_56_37 = g_56_41 | (p_56_41 & g_40_37);
 assign p_56_38 = p_56_41 & p_40_38;
 assign g_56_38 = g_56_41 | (p_56_41 & g_40_38);
 assign p_56_39 = p_56_41 & p_40_39;
 assign g_56_39 = g_56_41 | (p_56_41 & g_40_39);
 assign p_56_40 = p_56_41 & p_40_40;
 assign g_56_40 = g_56_41 | (p_56_41 & g_40_40);
 assign p_56_41 = p_56_49 & p_48_41;
 assign g_56_41 = g_56_49 | (p_56_49 & g_48_41);
 assign p_56_42 = p_56_49 & p_48_42;
 assign g_56_42 = g_56_49 | (p_56_49 & g_48_42);
 assign p_56_43 = p_56_49 & p_48_43;
 assign g_56_43 = g_56_49 | (p_56_49 & g_48_43);
 assign p_56_44 = p_56_49 & p_48_44;
 assign g_56_44 = g_56_49 | (p_56_49 & g_48_44);
 assign p_56_45 = p_56_49 & p_48_45;
 assign g_56_45 = g_56_49 | (p_56_49 & g_48_45);
 assign p_56_46 = p_56_49 & p_48_46;
 assign g_56_46 = g_56_49 | (p_56_49 & g_48_46);
 assign p_56_47 = p_56_49 & p_48_47;
 assign g_56_47 = g_56_49 | (p_56_49 & g_48_47);
 assign p_56_48 = p_56_49 & p_48_48;
 assign g_56_48 = g_56_49 | (p_56_49 & g_48_48);
 assign p_56_49 = p_56_53 & p_52_49;
 assign g_56_49 = g_56_53 | (p_56_53 & g_52_49);
 assign p_56_50 = p_56_53 & p_52_50;
 assign g_56_50 = g_56_53 | (p_56_53 & g_52_50);
 assign p_56_51 = p_56_53 & p_52_51;
 assign g_56_51 = g_56_53 | (p_56_53 & g_52_51);
 assign p_56_52 = p_56_53 & p_52_52;
 assign g_56_52 = g_56_53 | (p_56_53 & g_52_52);
 assign p_56_53 = p_56_55 & p_54_53;
 assign g_56_53 = g_56_55 | (p_56_55 & g_54_53);
 assign p_56_54 = p_56_55 & p_54_54;
 assign g_56_54 = g_56_55 | (p_56_55 & g_54_54);
 assign p_56_55 = p_56_56 & p_55_55;
 assign g_56_55 = g_56_56 | (p_56_56 & g_55_55);
 assign sum[56] = p_56_56^ g_55_0;
 assign p_57_0 = p_57_26 & p_25_0;
 assign g_57_0 = g_57_26 | (p_57_26 & g_25_0);
 assign p_57_1 = p_57_26 & p_25_1;
 assign g_57_1 = g_57_26 | (p_57_26 & g_25_1);
 assign p_57_2 = p_57_26 & p_25_2;
 assign g_57_2 = g_57_26 | (p_57_26 & g_25_2);
 assign p_57_3 = p_57_26 & p_25_3;
 assign g_57_3 = g_57_26 | (p_57_26 & g_25_3);
 assign p_57_4 = p_57_26 & p_25_4;
 assign g_57_4 = g_57_26 | (p_57_26 & g_25_4);
 assign p_57_5 = p_57_26 & p_25_5;
 assign g_57_5 = g_57_26 | (p_57_26 & g_25_5);
 assign p_57_6 = p_57_26 & p_25_6;
 assign g_57_6 = g_57_26 | (p_57_26 & g_25_6);
 assign p_57_7 = p_57_26 & p_25_7;
 assign g_57_7 = g_57_26 | (p_57_26 & g_25_7);
 assign p_57_8 = p_57_26 & p_25_8;
 assign g_57_8 = g_57_26 | (p_57_26 & g_25_8);
 assign p_57_9 = p_57_26 & p_25_9;
 assign g_57_9 = g_57_26 | (p_57_26 & g_25_9);
 assign p_57_10 = p_57_26 & p_25_10;
 assign g_57_10 = g_57_26 | (p_57_26 & g_25_10);
 assign p_57_11 = p_57_26 & p_25_11;
 assign g_57_11 = g_57_26 | (p_57_26 & g_25_11);
 assign p_57_12 = p_57_26 & p_25_12;
 assign g_57_12 = g_57_26 | (p_57_26 & g_25_12);
 assign p_57_13 = p_57_26 & p_25_13;
 assign g_57_13 = g_57_26 | (p_57_26 & g_25_13);
 assign p_57_14 = p_57_26 & p_25_14;
 assign g_57_14 = g_57_26 | (p_57_26 & g_25_14);
 assign p_57_15 = p_57_26 & p_25_15;
 assign g_57_15 = g_57_26 | (p_57_26 & g_25_15);
 assign p_57_16 = p_57_26 & p_25_16;
 assign g_57_16 = g_57_26 | (p_57_26 & g_25_16);
 assign p_57_17 = p_57_26 & p_25_17;
 assign g_57_17 = g_57_26 | (p_57_26 & g_25_17);
 assign p_57_18 = p_57_26 & p_25_18;
 assign g_57_18 = g_57_26 | (p_57_26 & g_25_18);
 assign p_57_19 = p_57_26 & p_25_19;
 assign g_57_19 = g_57_26 | (p_57_26 & g_25_19);
 assign p_57_20 = p_57_26 & p_25_20;
 assign g_57_20 = g_57_26 | (p_57_26 & g_25_20);
 assign p_57_21 = p_57_26 & p_25_21;
 assign g_57_21 = g_57_26 | (p_57_26 & g_25_21);
 assign p_57_22 = p_57_26 & p_25_22;
 assign g_57_22 = g_57_26 | (p_57_26 & g_25_22);
 assign p_57_23 = p_57_26 & p_25_23;
 assign g_57_23 = g_57_26 | (p_57_26 & g_25_23);
 assign p_57_24 = p_57_26 & p_25_24;
 assign g_57_24 = g_57_26 | (p_57_26 & g_25_24);
 assign p_57_25 = p_57_26 & p_25_25;
 assign g_57_25 = g_57_26 | (p_57_26 & g_25_25);
 assign p_57_26 = p_57_42 & p_41_26;
 assign g_57_26 = g_57_42 | (p_57_42 & g_41_26);
 assign p_57_27 = p_57_42 & p_41_27;
 assign g_57_27 = g_57_42 | (p_57_42 & g_41_27);
 assign p_57_28 = p_57_42 & p_41_28;
 assign g_57_28 = g_57_42 | (p_57_42 & g_41_28);
 assign p_57_29 = p_57_42 & p_41_29;
 assign g_57_29 = g_57_42 | (p_57_42 & g_41_29);
 assign p_57_30 = p_57_42 & p_41_30;
 assign g_57_30 = g_57_42 | (p_57_42 & g_41_30);
 assign p_57_31 = p_57_42 & p_41_31;
 assign g_57_31 = g_57_42 | (p_57_42 & g_41_31);
 assign p_57_32 = p_57_42 & p_41_32;
 assign g_57_32 = g_57_42 | (p_57_42 & g_41_32);
 assign p_57_33 = p_57_42 & p_41_33;
 assign g_57_33 = g_57_42 | (p_57_42 & g_41_33);
 assign p_57_34 = p_57_42 & p_41_34;
 assign g_57_34 = g_57_42 | (p_57_42 & g_41_34);
 assign p_57_35 = p_57_42 & p_41_35;
 assign g_57_35 = g_57_42 | (p_57_42 & g_41_35);
 assign p_57_36 = p_57_42 & p_41_36;
 assign g_57_36 = g_57_42 | (p_57_42 & g_41_36);
 assign p_57_37 = p_57_42 & p_41_37;
 assign g_57_37 = g_57_42 | (p_57_42 & g_41_37);
 assign p_57_38 = p_57_42 & p_41_38;
 assign g_57_38 = g_57_42 | (p_57_42 & g_41_38);
 assign p_57_39 = p_57_42 & p_41_39;
 assign g_57_39 = g_57_42 | (p_57_42 & g_41_39);
 assign p_57_40 = p_57_42 & p_41_40;
 assign g_57_40 = g_57_42 | (p_57_42 & g_41_40);
 assign p_57_41 = p_57_42 & p_41_41;
 assign g_57_41 = g_57_42 | (p_57_42 & g_41_41);
 assign p_57_42 = p_57_50 & p_49_42;
 assign g_57_42 = g_57_50 | (p_57_50 & g_49_42);
 assign p_57_43 = p_57_50 & p_49_43;
 assign g_57_43 = g_57_50 | (p_57_50 & g_49_43);
 assign p_57_44 = p_57_50 & p_49_44;
 assign g_57_44 = g_57_50 | (p_57_50 & g_49_44);
 assign p_57_45 = p_57_50 & p_49_45;
 assign g_57_45 = g_57_50 | (p_57_50 & g_49_45);
 assign p_57_46 = p_57_50 & p_49_46;
 assign g_57_46 = g_57_50 | (p_57_50 & g_49_46);
 assign p_57_47 = p_57_50 & p_49_47;
 assign g_57_47 = g_57_50 | (p_57_50 & g_49_47);
 assign p_57_48 = p_57_50 & p_49_48;
 assign g_57_48 = g_57_50 | (p_57_50 & g_49_48);
 assign p_57_49 = p_57_50 & p_49_49;
 assign g_57_49 = g_57_50 | (p_57_50 & g_49_49);
 assign p_57_50 = p_57_54 & p_53_50;
 assign g_57_50 = g_57_54 | (p_57_54 & g_53_50);
 assign p_57_51 = p_57_54 & p_53_51;
 assign g_57_51 = g_57_54 | (p_57_54 & g_53_51);
 assign p_57_52 = p_57_54 & p_53_52;
 assign g_57_52 = g_57_54 | (p_57_54 & g_53_52);
 assign p_57_53 = p_57_54 & p_53_53;
 assign g_57_53 = g_57_54 | (p_57_54 & g_53_53);
 assign p_57_54 = p_57_56 & p_55_54;
 assign g_57_54 = g_57_56 | (p_57_56 & g_55_54);
 assign p_57_55 = p_57_56 & p_55_55;
 assign g_57_55 = g_57_56 | (p_57_56 & g_55_55);
 assign p_57_56 = p_57_57 & p_56_56;
 assign g_57_56 = g_57_57 | (p_57_57 & g_56_56);
 assign sum[57] = p_57_57^ g_56_0;
 assign p_58_0 = p_58_27 & p_26_0;
 assign g_58_0 = g_58_27 | (p_58_27 & g_26_0);
 assign p_58_1 = p_58_27 & p_26_1;
 assign g_58_1 = g_58_27 | (p_58_27 & g_26_1);
 assign p_58_2 = p_58_27 & p_26_2;
 assign g_58_2 = g_58_27 | (p_58_27 & g_26_2);
 assign p_58_3 = p_58_27 & p_26_3;
 assign g_58_3 = g_58_27 | (p_58_27 & g_26_3);
 assign p_58_4 = p_58_27 & p_26_4;
 assign g_58_4 = g_58_27 | (p_58_27 & g_26_4);
 assign p_58_5 = p_58_27 & p_26_5;
 assign g_58_5 = g_58_27 | (p_58_27 & g_26_5);
 assign p_58_6 = p_58_27 & p_26_6;
 assign g_58_6 = g_58_27 | (p_58_27 & g_26_6);
 assign p_58_7 = p_58_27 & p_26_7;
 assign g_58_7 = g_58_27 | (p_58_27 & g_26_7);
 assign p_58_8 = p_58_27 & p_26_8;
 assign g_58_8 = g_58_27 | (p_58_27 & g_26_8);
 assign p_58_9 = p_58_27 & p_26_9;
 assign g_58_9 = g_58_27 | (p_58_27 & g_26_9);
 assign p_58_10 = p_58_27 & p_26_10;
 assign g_58_10 = g_58_27 | (p_58_27 & g_26_10);
 assign p_58_11 = p_58_27 & p_26_11;
 assign g_58_11 = g_58_27 | (p_58_27 & g_26_11);
 assign p_58_12 = p_58_27 & p_26_12;
 assign g_58_12 = g_58_27 | (p_58_27 & g_26_12);
 assign p_58_13 = p_58_27 & p_26_13;
 assign g_58_13 = g_58_27 | (p_58_27 & g_26_13);
 assign p_58_14 = p_58_27 & p_26_14;
 assign g_58_14 = g_58_27 | (p_58_27 & g_26_14);
 assign p_58_15 = p_58_27 & p_26_15;
 assign g_58_15 = g_58_27 | (p_58_27 & g_26_15);
 assign p_58_16 = p_58_27 & p_26_16;
 assign g_58_16 = g_58_27 | (p_58_27 & g_26_16);
 assign p_58_17 = p_58_27 & p_26_17;
 assign g_58_17 = g_58_27 | (p_58_27 & g_26_17);
 assign p_58_18 = p_58_27 & p_26_18;
 assign g_58_18 = g_58_27 | (p_58_27 & g_26_18);
 assign p_58_19 = p_58_27 & p_26_19;
 assign g_58_19 = g_58_27 | (p_58_27 & g_26_19);
 assign p_58_20 = p_58_27 & p_26_20;
 assign g_58_20 = g_58_27 | (p_58_27 & g_26_20);
 assign p_58_21 = p_58_27 & p_26_21;
 assign g_58_21 = g_58_27 | (p_58_27 & g_26_21);
 assign p_58_22 = p_58_27 & p_26_22;
 assign g_58_22 = g_58_27 | (p_58_27 & g_26_22);
 assign p_58_23 = p_58_27 & p_26_23;
 assign g_58_23 = g_58_27 | (p_58_27 & g_26_23);
 assign p_58_24 = p_58_27 & p_26_24;
 assign g_58_24 = g_58_27 | (p_58_27 & g_26_24);
 assign p_58_25 = p_58_27 & p_26_25;
 assign g_58_25 = g_58_27 | (p_58_27 & g_26_25);
 assign p_58_26 = p_58_27 & p_26_26;
 assign g_58_26 = g_58_27 | (p_58_27 & g_26_26);
 assign p_58_27 = p_58_43 & p_42_27;
 assign g_58_27 = g_58_43 | (p_58_43 & g_42_27);
 assign p_58_28 = p_58_43 & p_42_28;
 assign g_58_28 = g_58_43 | (p_58_43 & g_42_28);
 assign p_58_29 = p_58_43 & p_42_29;
 assign g_58_29 = g_58_43 | (p_58_43 & g_42_29);
 assign p_58_30 = p_58_43 & p_42_30;
 assign g_58_30 = g_58_43 | (p_58_43 & g_42_30);
 assign p_58_31 = p_58_43 & p_42_31;
 assign g_58_31 = g_58_43 | (p_58_43 & g_42_31);
 assign p_58_32 = p_58_43 & p_42_32;
 assign g_58_32 = g_58_43 | (p_58_43 & g_42_32);
 assign p_58_33 = p_58_43 & p_42_33;
 assign g_58_33 = g_58_43 | (p_58_43 & g_42_33);
 assign p_58_34 = p_58_43 & p_42_34;
 assign g_58_34 = g_58_43 | (p_58_43 & g_42_34);
 assign p_58_35 = p_58_43 & p_42_35;
 assign g_58_35 = g_58_43 | (p_58_43 & g_42_35);
 assign p_58_36 = p_58_43 & p_42_36;
 assign g_58_36 = g_58_43 | (p_58_43 & g_42_36);
 assign p_58_37 = p_58_43 & p_42_37;
 assign g_58_37 = g_58_43 | (p_58_43 & g_42_37);
 assign p_58_38 = p_58_43 & p_42_38;
 assign g_58_38 = g_58_43 | (p_58_43 & g_42_38);
 assign p_58_39 = p_58_43 & p_42_39;
 assign g_58_39 = g_58_43 | (p_58_43 & g_42_39);
 assign p_58_40 = p_58_43 & p_42_40;
 assign g_58_40 = g_58_43 | (p_58_43 & g_42_40);
 assign p_58_41 = p_58_43 & p_42_41;
 assign g_58_41 = g_58_43 | (p_58_43 & g_42_41);
 assign p_58_42 = p_58_43 & p_42_42;
 assign g_58_42 = g_58_43 | (p_58_43 & g_42_42);
 assign p_58_43 = p_58_51 & p_50_43;
 assign g_58_43 = g_58_51 | (p_58_51 & g_50_43);
 assign p_58_44 = p_58_51 & p_50_44;
 assign g_58_44 = g_58_51 | (p_58_51 & g_50_44);
 assign p_58_45 = p_58_51 & p_50_45;
 assign g_58_45 = g_58_51 | (p_58_51 & g_50_45);
 assign p_58_46 = p_58_51 & p_50_46;
 assign g_58_46 = g_58_51 | (p_58_51 & g_50_46);
 assign p_58_47 = p_58_51 & p_50_47;
 assign g_58_47 = g_58_51 | (p_58_51 & g_50_47);
 assign p_58_48 = p_58_51 & p_50_48;
 assign g_58_48 = g_58_51 | (p_58_51 & g_50_48);
 assign p_58_49 = p_58_51 & p_50_49;
 assign g_58_49 = g_58_51 | (p_58_51 & g_50_49);
 assign p_58_50 = p_58_51 & p_50_50;
 assign g_58_50 = g_58_51 | (p_58_51 & g_50_50);
 assign p_58_51 = p_58_55 & p_54_51;
 assign g_58_51 = g_58_55 | (p_58_55 & g_54_51);
 assign p_58_52 = p_58_55 & p_54_52;
 assign g_58_52 = g_58_55 | (p_58_55 & g_54_52);
 assign p_58_53 = p_58_55 & p_54_53;
 assign g_58_53 = g_58_55 | (p_58_55 & g_54_53);
 assign p_58_54 = p_58_55 & p_54_54;
 assign g_58_54 = g_58_55 | (p_58_55 & g_54_54);
 assign p_58_55 = p_58_57 & p_56_55;
 assign g_58_55 = g_58_57 | (p_58_57 & g_56_55);
 assign p_58_56 = p_58_57 & p_56_56;
 assign g_58_56 = g_58_57 | (p_58_57 & g_56_56);
 assign p_58_57 = p_58_58 & p_57_57;
 assign g_58_57 = g_58_58 | (p_58_58 & g_57_57);
 assign sum[58] = p_58_58^ g_57_0;
 assign p_59_0 = p_59_28 & p_27_0;
 assign g_59_0 = g_59_28 | (p_59_28 & g_27_0);
 assign p_59_1 = p_59_28 & p_27_1;
 assign g_59_1 = g_59_28 | (p_59_28 & g_27_1);
 assign p_59_2 = p_59_28 & p_27_2;
 assign g_59_2 = g_59_28 | (p_59_28 & g_27_2);
 assign p_59_3 = p_59_28 & p_27_3;
 assign g_59_3 = g_59_28 | (p_59_28 & g_27_3);
 assign p_59_4 = p_59_28 & p_27_4;
 assign g_59_4 = g_59_28 | (p_59_28 & g_27_4);
 assign p_59_5 = p_59_28 & p_27_5;
 assign g_59_5 = g_59_28 | (p_59_28 & g_27_5);
 assign p_59_6 = p_59_28 & p_27_6;
 assign g_59_6 = g_59_28 | (p_59_28 & g_27_6);
 assign p_59_7 = p_59_28 & p_27_7;
 assign g_59_7 = g_59_28 | (p_59_28 & g_27_7);
 assign p_59_8 = p_59_28 & p_27_8;
 assign g_59_8 = g_59_28 | (p_59_28 & g_27_8);
 assign p_59_9 = p_59_28 & p_27_9;
 assign g_59_9 = g_59_28 | (p_59_28 & g_27_9);
 assign p_59_10 = p_59_28 & p_27_10;
 assign g_59_10 = g_59_28 | (p_59_28 & g_27_10);
 assign p_59_11 = p_59_28 & p_27_11;
 assign g_59_11 = g_59_28 | (p_59_28 & g_27_11);
 assign p_59_12 = p_59_28 & p_27_12;
 assign g_59_12 = g_59_28 | (p_59_28 & g_27_12);
 assign p_59_13 = p_59_28 & p_27_13;
 assign g_59_13 = g_59_28 | (p_59_28 & g_27_13);
 assign p_59_14 = p_59_28 & p_27_14;
 assign g_59_14 = g_59_28 | (p_59_28 & g_27_14);
 assign p_59_15 = p_59_28 & p_27_15;
 assign g_59_15 = g_59_28 | (p_59_28 & g_27_15);
 assign p_59_16 = p_59_28 & p_27_16;
 assign g_59_16 = g_59_28 | (p_59_28 & g_27_16);
 assign p_59_17 = p_59_28 & p_27_17;
 assign g_59_17 = g_59_28 | (p_59_28 & g_27_17);
 assign p_59_18 = p_59_28 & p_27_18;
 assign g_59_18 = g_59_28 | (p_59_28 & g_27_18);
 assign p_59_19 = p_59_28 & p_27_19;
 assign g_59_19 = g_59_28 | (p_59_28 & g_27_19);
 assign p_59_20 = p_59_28 & p_27_20;
 assign g_59_20 = g_59_28 | (p_59_28 & g_27_20);
 assign p_59_21 = p_59_28 & p_27_21;
 assign g_59_21 = g_59_28 | (p_59_28 & g_27_21);
 assign p_59_22 = p_59_28 & p_27_22;
 assign g_59_22 = g_59_28 | (p_59_28 & g_27_22);
 assign p_59_23 = p_59_28 & p_27_23;
 assign g_59_23 = g_59_28 | (p_59_28 & g_27_23);
 assign p_59_24 = p_59_28 & p_27_24;
 assign g_59_24 = g_59_28 | (p_59_28 & g_27_24);
 assign p_59_25 = p_59_28 & p_27_25;
 assign g_59_25 = g_59_28 | (p_59_28 & g_27_25);
 assign p_59_26 = p_59_28 & p_27_26;
 assign g_59_26 = g_59_28 | (p_59_28 & g_27_26);
 assign p_59_27 = p_59_28 & p_27_27;
 assign g_59_27 = g_59_28 | (p_59_28 & g_27_27);
 assign p_59_28 = p_59_44 & p_43_28;
 assign g_59_28 = g_59_44 | (p_59_44 & g_43_28);
 assign p_59_29 = p_59_44 & p_43_29;
 assign g_59_29 = g_59_44 | (p_59_44 & g_43_29);
 assign p_59_30 = p_59_44 & p_43_30;
 assign g_59_30 = g_59_44 | (p_59_44 & g_43_30);
 assign p_59_31 = p_59_44 & p_43_31;
 assign g_59_31 = g_59_44 | (p_59_44 & g_43_31);
 assign p_59_32 = p_59_44 & p_43_32;
 assign g_59_32 = g_59_44 | (p_59_44 & g_43_32);
 assign p_59_33 = p_59_44 & p_43_33;
 assign g_59_33 = g_59_44 | (p_59_44 & g_43_33);
 assign p_59_34 = p_59_44 & p_43_34;
 assign g_59_34 = g_59_44 | (p_59_44 & g_43_34);
 assign p_59_35 = p_59_44 & p_43_35;
 assign g_59_35 = g_59_44 | (p_59_44 & g_43_35);
 assign p_59_36 = p_59_44 & p_43_36;
 assign g_59_36 = g_59_44 | (p_59_44 & g_43_36);
 assign p_59_37 = p_59_44 & p_43_37;
 assign g_59_37 = g_59_44 | (p_59_44 & g_43_37);
 assign p_59_38 = p_59_44 & p_43_38;
 assign g_59_38 = g_59_44 | (p_59_44 & g_43_38);
 assign p_59_39 = p_59_44 & p_43_39;
 assign g_59_39 = g_59_44 | (p_59_44 & g_43_39);
 assign p_59_40 = p_59_44 & p_43_40;
 assign g_59_40 = g_59_44 | (p_59_44 & g_43_40);
 assign p_59_41 = p_59_44 & p_43_41;
 assign g_59_41 = g_59_44 | (p_59_44 & g_43_41);
 assign p_59_42 = p_59_44 & p_43_42;
 assign g_59_42 = g_59_44 | (p_59_44 & g_43_42);
 assign p_59_43 = p_59_44 & p_43_43;
 assign g_59_43 = g_59_44 | (p_59_44 & g_43_43);
 assign p_59_44 = p_59_52 & p_51_44;
 assign g_59_44 = g_59_52 | (p_59_52 & g_51_44);
 assign p_59_45 = p_59_52 & p_51_45;
 assign g_59_45 = g_59_52 | (p_59_52 & g_51_45);
 assign p_59_46 = p_59_52 & p_51_46;
 assign g_59_46 = g_59_52 | (p_59_52 & g_51_46);
 assign p_59_47 = p_59_52 & p_51_47;
 assign g_59_47 = g_59_52 | (p_59_52 & g_51_47);
 assign p_59_48 = p_59_52 & p_51_48;
 assign g_59_48 = g_59_52 | (p_59_52 & g_51_48);
 assign p_59_49 = p_59_52 & p_51_49;
 assign g_59_49 = g_59_52 | (p_59_52 & g_51_49);
 assign p_59_50 = p_59_52 & p_51_50;
 assign g_59_50 = g_59_52 | (p_59_52 & g_51_50);
 assign p_59_51 = p_59_52 & p_51_51;
 assign g_59_51 = g_59_52 | (p_59_52 & g_51_51);
 assign p_59_52 = p_59_56 & p_55_52;
 assign g_59_52 = g_59_56 | (p_59_56 & g_55_52);
 assign p_59_53 = p_59_56 & p_55_53;
 assign g_59_53 = g_59_56 | (p_59_56 & g_55_53);
 assign p_59_54 = p_59_56 & p_55_54;
 assign g_59_54 = g_59_56 | (p_59_56 & g_55_54);
 assign p_59_55 = p_59_56 & p_55_55;
 assign g_59_55 = g_59_56 | (p_59_56 & g_55_55);
 assign p_59_56 = p_59_58 & p_57_56;
 assign g_59_56 = g_59_58 | (p_59_58 & g_57_56);
 assign p_59_57 = p_59_58 & p_57_57;
 assign g_59_57 = g_59_58 | (p_59_58 & g_57_57);
 assign p_59_58 = p_59_59 & p_58_58;
 assign g_59_58 = g_59_59 | (p_59_59 & g_58_58);
 assign sum[59] = p_59_59^ g_58_0;
 assign p_60_0 = p_60_29 & p_28_0;
 assign g_60_0 = g_60_29 | (p_60_29 & g_28_0);
 assign p_60_1 = p_60_29 & p_28_1;
 assign g_60_1 = g_60_29 | (p_60_29 & g_28_1);
 assign p_60_2 = p_60_29 & p_28_2;
 assign g_60_2 = g_60_29 | (p_60_29 & g_28_2);
 assign p_60_3 = p_60_29 & p_28_3;
 assign g_60_3 = g_60_29 | (p_60_29 & g_28_3);
 assign p_60_4 = p_60_29 & p_28_4;
 assign g_60_4 = g_60_29 | (p_60_29 & g_28_4);
 assign p_60_5 = p_60_29 & p_28_5;
 assign g_60_5 = g_60_29 | (p_60_29 & g_28_5);
 assign p_60_6 = p_60_29 & p_28_6;
 assign g_60_6 = g_60_29 | (p_60_29 & g_28_6);
 assign p_60_7 = p_60_29 & p_28_7;
 assign g_60_7 = g_60_29 | (p_60_29 & g_28_7);
 assign p_60_8 = p_60_29 & p_28_8;
 assign g_60_8 = g_60_29 | (p_60_29 & g_28_8);
 assign p_60_9 = p_60_29 & p_28_9;
 assign g_60_9 = g_60_29 | (p_60_29 & g_28_9);
 assign p_60_10 = p_60_29 & p_28_10;
 assign g_60_10 = g_60_29 | (p_60_29 & g_28_10);
 assign p_60_11 = p_60_29 & p_28_11;
 assign g_60_11 = g_60_29 | (p_60_29 & g_28_11);
 assign p_60_12 = p_60_29 & p_28_12;
 assign g_60_12 = g_60_29 | (p_60_29 & g_28_12);
 assign p_60_13 = p_60_29 & p_28_13;
 assign g_60_13 = g_60_29 | (p_60_29 & g_28_13);
 assign p_60_14 = p_60_29 & p_28_14;
 assign g_60_14 = g_60_29 | (p_60_29 & g_28_14);
 assign p_60_15 = p_60_29 & p_28_15;
 assign g_60_15 = g_60_29 | (p_60_29 & g_28_15);
 assign p_60_16 = p_60_29 & p_28_16;
 assign g_60_16 = g_60_29 | (p_60_29 & g_28_16);
 assign p_60_17 = p_60_29 & p_28_17;
 assign g_60_17 = g_60_29 | (p_60_29 & g_28_17);
 assign p_60_18 = p_60_29 & p_28_18;
 assign g_60_18 = g_60_29 | (p_60_29 & g_28_18);
 assign p_60_19 = p_60_29 & p_28_19;
 assign g_60_19 = g_60_29 | (p_60_29 & g_28_19);
 assign p_60_20 = p_60_29 & p_28_20;
 assign g_60_20 = g_60_29 | (p_60_29 & g_28_20);
 assign p_60_21 = p_60_29 & p_28_21;
 assign g_60_21 = g_60_29 | (p_60_29 & g_28_21);
 assign p_60_22 = p_60_29 & p_28_22;
 assign g_60_22 = g_60_29 | (p_60_29 & g_28_22);
 assign p_60_23 = p_60_29 & p_28_23;
 assign g_60_23 = g_60_29 | (p_60_29 & g_28_23);
 assign p_60_24 = p_60_29 & p_28_24;
 assign g_60_24 = g_60_29 | (p_60_29 & g_28_24);
 assign p_60_25 = p_60_29 & p_28_25;
 assign g_60_25 = g_60_29 | (p_60_29 & g_28_25);
 assign p_60_26 = p_60_29 & p_28_26;
 assign g_60_26 = g_60_29 | (p_60_29 & g_28_26);
 assign p_60_27 = p_60_29 & p_28_27;
 assign g_60_27 = g_60_29 | (p_60_29 & g_28_27);
 assign p_60_28 = p_60_29 & p_28_28;
 assign g_60_28 = g_60_29 | (p_60_29 & g_28_28);
 assign p_60_29 = p_60_45 & p_44_29;
 assign g_60_29 = g_60_45 | (p_60_45 & g_44_29);
 assign p_60_30 = p_60_45 & p_44_30;
 assign g_60_30 = g_60_45 | (p_60_45 & g_44_30);
 assign p_60_31 = p_60_45 & p_44_31;
 assign g_60_31 = g_60_45 | (p_60_45 & g_44_31);
 assign p_60_32 = p_60_45 & p_44_32;
 assign g_60_32 = g_60_45 | (p_60_45 & g_44_32);
 assign p_60_33 = p_60_45 & p_44_33;
 assign g_60_33 = g_60_45 | (p_60_45 & g_44_33);
 assign p_60_34 = p_60_45 & p_44_34;
 assign g_60_34 = g_60_45 | (p_60_45 & g_44_34);
 assign p_60_35 = p_60_45 & p_44_35;
 assign g_60_35 = g_60_45 | (p_60_45 & g_44_35);
 assign p_60_36 = p_60_45 & p_44_36;
 assign g_60_36 = g_60_45 | (p_60_45 & g_44_36);
 assign p_60_37 = p_60_45 & p_44_37;
 assign g_60_37 = g_60_45 | (p_60_45 & g_44_37);
 assign p_60_38 = p_60_45 & p_44_38;
 assign g_60_38 = g_60_45 | (p_60_45 & g_44_38);
 assign p_60_39 = p_60_45 & p_44_39;
 assign g_60_39 = g_60_45 | (p_60_45 & g_44_39);
 assign p_60_40 = p_60_45 & p_44_40;
 assign g_60_40 = g_60_45 | (p_60_45 & g_44_40);
 assign p_60_41 = p_60_45 & p_44_41;
 assign g_60_41 = g_60_45 | (p_60_45 & g_44_41);
 assign p_60_42 = p_60_45 & p_44_42;
 assign g_60_42 = g_60_45 | (p_60_45 & g_44_42);
 assign p_60_43 = p_60_45 & p_44_43;
 assign g_60_43 = g_60_45 | (p_60_45 & g_44_43);
 assign p_60_44 = p_60_45 & p_44_44;
 assign g_60_44 = g_60_45 | (p_60_45 & g_44_44);
 assign p_60_45 = p_60_53 & p_52_45;
 assign g_60_45 = g_60_53 | (p_60_53 & g_52_45);
 assign p_60_46 = p_60_53 & p_52_46;
 assign g_60_46 = g_60_53 | (p_60_53 & g_52_46);
 assign p_60_47 = p_60_53 & p_52_47;
 assign g_60_47 = g_60_53 | (p_60_53 & g_52_47);
 assign p_60_48 = p_60_53 & p_52_48;
 assign g_60_48 = g_60_53 | (p_60_53 & g_52_48);
 assign p_60_49 = p_60_53 & p_52_49;
 assign g_60_49 = g_60_53 | (p_60_53 & g_52_49);
 assign p_60_50 = p_60_53 & p_52_50;
 assign g_60_50 = g_60_53 | (p_60_53 & g_52_50);
 assign p_60_51 = p_60_53 & p_52_51;
 assign g_60_51 = g_60_53 | (p_60_53 & g_52_51);
 assign p_60_52 = p_60_53 & p_52_52;
 assign g_60_52 = g_60_53 | (p_60_53 & g_52_52);
 assign p_60_53 = p_60_57 & p_56_53;
 assign g_60_53 = g_60_57 | (p_60_57 & g_56_53);
 assign p_60_54 = p_60_57 & p_56_54;
 assign g_60_54 = g_60_57 | (p_60_57 & g_56_54);
 assign p_60_55 = p_60_57 & p_56_55;
 assign g_60_55 = g_60_57 | (p_60_57 & g_56_55);
 assign p_60_56 = p_60_57 & p_56_56;
 assign g_60_56 = g_60_57 | (p_60_57 & g_56_56);
 assign p_60_57 = p_60_59 & p_58_57;
 assign g_60_57 = g_60_59 | (p_60_59 & g_58_57);
 assign p_60_58 = p_60_59 & p_58_58;
 assign g_60_58 = g_60_59 | (p_60_59 & g_58_58);
 assign p_60_59 = p_60_60 & p_59_59;
 assign g_60_59 = g_60_60 | (p_60_60 & g_59_59);
 assign sum[60] = p_60_60^ g_59_0;
 assign p_61_0 = p_61_30 & p_29_0;
 assign g_61_0 = g_61_30 | (p_61_30 & g_29_0);
 assign p_61_1 = p_61_30 & p_29_1;
 assign g_61_1 = g_61_30 | (p_61_30 & g_29_1);
 assign p_61_2 = p_61_30 & p_29_2;
 assign g_61_2 = g_61_30 | (p_61_30 & g_29_2);
 assign p_61_3 = p_61_30 & p_29_3;
 assign g_61_3 = g_61_30 | (p_61_30 & g_29_3);
 assign p_61_4 = p_61_30 & p_29_4;
 assign g_61_4 = g_61_30 | (p_61_30 & g_29_4);
 assign p_61_5 = p_61_30 & p_29_5;
 assign g_61_5 = g_61_30 | (p_61_30 & g_29_5);
 assign p_61_6 = p_61_30 & p_29_6;
 assign g_61_6 = g_61_30 | (p_61_30 & g_29_6);
 assign p_61_7 = p_61_30 & p_29_7;
 assign g_61_7 = g_61_30 | (p_61_30 & g_29_7);
 assign p_61_8 = p_61_30 & p_29_8;
 assign g_61_8 = g_61_30 | (p_61_30 & g_29_8);
 assign p_61_9 = p_61_30 & p_29_9;
 assign g_61_9 = g_61_30 | (p_61_30 & g_29_9);
 assign p_61_10 = p_61_30 & p_29_10;
 assign g_61_10 = g_61_30 | (p_61_30 & g_29_10);
 assign p_61_11 = p_61_30 & p_29_11;
 assign g_61_11 = g_61_30 | (p_61_30 & g_29_11);
 assign p_61_12 = p_61_30 & p_29_12;
 assign g_61_12 = g_61_30 | (p_61_30 & g_29_12);
 assign p_61_13 = p_61_30 & p_29_13;
 assign g_61_13 = g_61_30 | (p_61_30 & g_29_13);
 assign p_61_14 = p_61_30 & p_29_14;
 assign g_61_14 = g_61_30 | (p_61_30 & g_29_14);
 assign p_61_15 = p_61_30 & p_29_15;
 assign g_61_15 = g_61_30 | (p_61_30 & g_29_15);
 assign p_61_16 = p_61_30 & p_29_16;
 assign g_61_16 = g_61_30 | (p_61_30 & g_29_16);
 assign p_61_17 = p_61_30 & p_29_17;
 assign g_61_17 = g_61_30 | (p_61_30 & g_29_17);
 assign p_61_18 = p_61_30 & p_29_18;
 assign g_61_18 = g_61_30 | (p_61_30 & g_29_18);
 assign p_61_19 = p_61_30 & p_29_19;
 assign g_61_19 = g_61_30 | (p_61_30 & g_29_19);
 assign p_61_20 = p_61_30 & p_29_20;
 assign g_61_20 = g_61_30 | (p_61_30 & g_29_20);
 assign p_61_21 = p_61_30 & p_29_21;
 assign g_61_21 = g_61_30 | (p_61_30 & g_29_21);
 assign p_61_22 = p_61_30 & p_29_22;
 assign g_61_22 = g_61_30 | (p_61_30 & g_29_22);
 assign p_61_23 = p_61_30 & p_29_23;
 assign g_61_23 = g_61_30 | (p_61_30 & g_29_23);
 assign p_61_24 = p_61_30 & p_29_24;
 assign g_61_24 = g_61_30 | (p_61_30 & g_29_24);
 assign p_61_25 = p_61_30 & p_29_25;
 assign g_61_25 = g_61_30 | (p_61_30 & g_29_25);
 assign p_61_26 = p_61_30 & p_29_26;
 assign g_61_26 = g_61_30 | (p_61_30 & g_29_26);
 assign p_61_27 = p_61_30 & p_29_27;
 assign g_61_27 = g_61_30 | (p_61_30 & g_29_27);
 assign p_61_28 = p_61_30 & p_29_28;
 assign g_61_28 = g_61_30 | (p_61_30 & g_29_28);
 assign p_61_29 = p_61_30 & p_29_29;
 assign g_61_29 = g_61_30 | (p_61_30 & g_29_29);
 assign p_61_30 = p_61_46 & p_45_30;
 assign g_61_30 = g_61_46 | (p_61_46 & g_45_30);
 assign p_61_31 = p_61_46 & p_45_31;
 assign g_61_31 = g_61_46 | (p_61_46 & g_45_31);
 assign p_61_32 = p_61_46 & p_45_32;
 assign g_61_32 = g_61_46 | (p_61_46 & g_45_32);
 assign p_61_33 = p_61_46 & p_45_33;
 assign g_61_33 = g_61_46 | (p_61_46 & g_45_33);
 assign p_61_34 = p_61_46 & p_45_34;
 assign g_61_34 = g_61_46 | (p_61_46 & g_45_34);
 assign p_61_35 = p_61_46 & p_45_35;
 assign g_61_35 = g_61_46 | (p_61_46 & g_45_35);
 assign p_61_36 = p_61_46 & p_45_36;
 assign g_61_36 = g_61_46 | (p_61_46 & g_45_36);
 assign p_61_37 = p_61_46 & p_45_37;
 assign g_61_37 = g_61_46 | (p_61_46 & g_45_37);
 assign p_61_38 = p_61_46 & p_45_38;
 assign g_61_38 = g_61_46 | (p_61_46 & g_45_38);
 assign p_61_39 = p_61_46 & p_45_39;
 assign g_61_39 = g_61_46 | (p_61_46 & g_45_39);
 assign p_61_40 = p_61_46 & p_45_40;
 assign g_61_40 = g_61_46 | (p_61_46 & g_45_40);
 assign p_61_41 = p_61_46 & p_45_41;
 assign g_61_41 = g_61_46 | (p_61_46 & g_45_41);
 assign p_61_42 = p_61_46 & p_45_42;
 assign g_61_42 = g_61_46 | (p_61_46 & g_45_42);
 assign p_61_43 = p_61_46 & p_45_43;
 assign g_61_43 = g_61_46 | (p_61_46 & g_45_43);
 assign p_61_44 = p_61_46 & p_45_44;
 assign g_61_44 = g_61_46 | (p_61_46 & g_45_44);
 assign p_61_45 = p_61_46 & p_45_45;
 assign g_61_45 = g_61_46 | (p_61_46 & g_45_45);
 assign p_61_46 = p_61_54 & p_53_46;
 assign g_61_46 = g_61_54 | (p_61_54 & g_53_46);
 assign p_61_47 = p_61_54 & p_53_47;
 assign g_61_47 = g_61_54 | (p_61_54 & g_53_47);
 assign p_61_48 = p_61_54 & p_53_48;
 assign g_61_48 = g_61_54 | (p_61_54 & g_53_48);
 assign p_61_49 = p_61_54 & p_53_49;
 assign g_61_49 = g_61_54 | (p_61_54 & g_53_49);
 assign p_61_50 = p_61_54 & p_53_50;
 assign g_61_50 = g_61_54 | (p_61_54 & g_53_50);
 assign p_61_51 = p_61_54 & p_53_51;
 assign g_61_51 = g_61_54 | (p_61_54 & g_53_51);
 assign p_61_52 = p_61_54 & p_53_52;
 assign g_61_52 = g_61_54 | (p_61_54 & g_53_52);
 assign p_61_53 = p_61_54 & p_53_53;
 assign g_61_53 = g_61_54 | (p_61_54 & g_53_53);
 assign p_61_54 = p_61_58 & p_57_54;
 assign g_61_54 = g_61_58 | (p_61_58 & g_57_54);
 assign p_61_55 = p_61_58 & p_57_55;
 assign g_61_55 = g_61_58 | (p_61_58 & g_57_55);
 assign p_61_56 = p_61_58 & p_57_56;
 assign g_61_56 = g_61_58 | (p_61_58 & g_57_56);
 assign p_61_57 = p_61_58 & p_57_57;
 assign g_61_57 = g_61_58 | (p_61_58 & g_57_57);
 assign p_61_58 = p_61_60 & p_59_58;
 assign g_61_58 = g_61_60 | (p_61_60 & g_59_58);
 assign p_61_59 = p_61_60 & p_59_59;
 assign g_61_59 = g_61_60 | (p_61_60 & g_59_59);
 assign p_61_60 = p_61_61 & p_60_60;
 assign g_61_60 = g_61_61 | (p_61_61 & g_60_60);
 assign sum[61] = p_61_61^ g_60_0;
 assign p_62_0 = p_62_31 & p_30_0;
 assign g_62_0 = g_62_31 | (p_62_31 & g_30_0);
 assign p_62_1 = p_62_31 & p_30_1;
 assign g_62_1 = g_62_31 | (p_62_31 & g_30_1);
 assign p_62_2 = p_62_31 & p_30_2;
 assign g_62_2 = g_62_31 | (p_62_31 & g_30_2);
 assign p_62_3 = p_62_31 & p_30_3;
 assign g_62_3 = g_62_31 | (p_62_31 & g_30_3);
 assign p_62_4 = p_62_31 & p_30_4;
 assign g_62_4 = g_62_31 | (p_62_31 & g_30_4);
 assign p_62_5 = p_62_31 & p_30_5;
 assign g_62_5 = g_62_31 | (p_62_31 & g_30_5);
 assign p_62_6 = p_62_31 & p_30_6;
 assign g_62_6 = g_62_31 | (p_62_31 & g_30_6);
 assign p_62_7 = p_62_31 & p_30_7;
 assign g_62_7 = g_62_31 | (p_62_31 & g_30_7);
 assign p_62_8 = p_62_31 & p_30_8;
 assign g_62_8 = g_62_31 | (p_62_31 & g_30_8);
 assign p_62_9 = p_62_31 & p_30_9;
 assign g_62_9 = g_62_31 | (p_62_31 & g_30_9);
 assign p_62_10 = p_62_31 & p_30_10;
 assign g_62_10 = g_62_31 | (p_62_31 & g_30_10);
 assign p_62_11 = p_62_31 & p_30_11;
 assign g_62_11 = g_62_31 | (p_62_31 & g_30_11);
 assign p_62_12 = p_62_31 & p_30_12;
 assign g_62_12 = g_62_31 | (p_62_31 & g_30_12);
 assign p_62_13 = p_62_31 & p_30_13;
 assign g_62_13 = g_62_31 | (p_62_31 & g_30_13);
 assign p_62_14 = p_62_31 & p_30_14;
 assign g_62_14 = g_62_31 | (p_62_31 & g_30_14);
 assign p_62_15 = p_62_31 & p_30_15;
 assign g_62_15 = g_62_31 | (p_62_31 & g_30_15);
 assign p_62_16 = p_62_31 & p_30_16;
 assign g_62_16 = g_62_31 | (p_62_31 & g_30_16);
 assign p_62_17 = p_62_31 & p_30_17;
 assign g_62_17 = g_62_31 | (p_62_31 & g_30_17);
 assign p_62_18 = p_62_31 & p_30_18;
 assign g_62_18 = g_62_31 | (p_62_31 & g_30_18);
 assign p_62_19 = p_62_31 & p_30_19;
 assign g_62_19 = g_62_31 | (p_62_31 & g_30_19);
 assign p_62_20 = p_62_31 & p_30_20;
 assign g_62_20 = g_62_31 | (p_62_31 & g_30_20);
 assign p_62_21 = p_62_31 & p_30_21;
 assign g_62_21 = g_62_31 | (p_62_31 & g_30_21);
 assign p_62_22 = p_62_31 & p_30_22;
 assign g_62_22 = g_62_31 | (p_62_31 & g_30_22);
 assign p_62_23 = p_62_31 & p_30_23;
 assign g_62_23 = g_62_31 | (p_62_31 & g_30_23);
 assign p_62_24 = p_62_31 & p_30_24;
 assign g_62_24 = g_62_31 | (p_62_31 & g_30_24);
 assign p_62_25 = p_62_31 & p_30_25;
 assign g_62_25 = g_62_31 | (p_62_31 & g_30_25);
 assign p_62_26 = p_62_31 & p_30_26;
 assign g_62_26 = g_62_31 | (p_62_31 & g_30_26);
 assign p_62_27 = p_62_31 & p_30_27;
 assign g_62_27 = g_62_31 | (p_62_31 & g_30_27);
 assign p_62_28 = p_62_31 & p_30_28;
 assign g_62_28 = g_62_31 | (p_62_31 & g_30_28);
 assign p_62_29 = p_62_31 & p_30_29;
 assign g_62_29 = g_62_31 | (p_62_31 & g_30_29);
 assign p_62_30 = p_62_31 & p_30_30;
 assign g_62_30 = g_62_31 | (p_62_31 & g_30_30);
 assign p_62_31 = p_62_47 & p_46_31;
 assign g_62_31 = g_62_47 | (p_62_47 & g_46_31);
 assign p_62_32 = p_62_47 & p_46_32;
 assign g_62_32 = g_62_47 | (p_62_47 & g_46_32);
 assign p_62_33 = p_62_47 & p_46_33;
 assign g_62_33 = g_62_47 | (p_62_47 & g_46_33);
 assign p_62_34 = p_62_47 & p_46_34;
 assign g_62_34 = g_62_47 | (p_62_47 & g_46_34);
 assign p_62_35 = p_62_47 & p_46_35;
 assign g_62_35 = g_62_47 | (p_62_47 & g_46_35);
 assign p_62_36 = p_62_47 & p_46_36;
 assign g_62_36 = g_62_47 | (p_62_47 & g_46_36);
 assign p_62_37 = p_62_47 & p_46_37;
 assign g_62_37 = g_62_47 | (p_62_47 & g_46_37);
 assign p_62_38 = p_62_47 & p_46_38;
 assign g_62_38 = g_62_47 | (p_62_47 & g_46_38);
 assign p_62_39 = p_62_47 & p_46_39;
 assign g_62_39 = g_62_47 | (p_62_47 & g_46_39);
 assign p_62_40 = p_62_47 & p_46_40;
 assign g_62_40 = g_62_47 | (p_62_47 & g_46_40);
 assign p_62_41 = p_62_47 & p_46_41;
 assign g_62_41 = g_62_47 | (p_62_47 & g_46_41);
 assign p_62_42 = p_62_47 & p_46_42;
 assign g_62_42 = g_62_47 | (p_62_47 & g_46_42);
 assign p_62_43 = p_62_47 & p_46_43;
 assign g_62_43 = g_62_47 | (p_62_47 & g_46_43);
 assign p_62_44 = p_62_47 & p_46_44;
 assign g_62_44 = g_62_47 | (p_62_47 & g_46_44);
 assign p_62_45 = p_62_47 & p_46_45;
 assign g_62_45 = g_62_47 | (p_62_47 & g_46_45);
 assign p_62_46 = p_62_47 & p_46_46;
 assign g_62_46 = g_62_47 | (p_62_47 & g_46_46);
 assign p_62_47 = p_62_55 & p_54_47;
 assign g_62_47 = g_62_55 | (p_62_55 & g_54_47);
 assign p_62_48 = p_62_55 & p_54_48;
 assign g_62_48 = g_62_55 | (p_62_55 & g_54_48);
 assign p_62_49 = p_62_55 & p_54_49;
 assign g_62_49 = g_62_55 | (p_62_55 & g_54_49);
 assign p_62_50 = p_62_55 & p_54_50;
 assign g_62_50 = g_62_55 | (p_62_55 & g_54_50);
 assign p_62_51 = p_62_55 & p_54_51;
 assign g_62_51 = g_62_55 | (p_62_55 & g_54_51);
 assign p_62_52 = p_62_55 & p_54_52;
 assign g_62_52 = g_62_55 | (p_62_55 & g_54_52);
 assign p_62_53 = p_62_55 & p_54_53;
 assign g_62_53 = g_62_55 | (p_62_55 & g_54_53);
 assign p_62_54 = p_62_55 & p_54_54;
 assign g_62_54 = g_62_55 | (p_62_55 & g_54_54);
 assign p_62_55 = p_62_59 & p_58_55;
 assign g_62_55 = g_62_59 | (p_62_59 & g_58_55);
 assign p_62_56 = p_62_59 & p_58_56;
 assign g_62_56 = g_62_59 | (p_62_59 & g_58_56);
 assign p_62_57 = p_62_59 & p_58_57;
 assign g_62_57 = g_62_59 | (p_62_59 & g_58_57);
 assign p_62_58 = p_62_59 & p_58_58;
 assign g_62_58 = g_62_59 | (p_62_59 & g_58_58);
 assign p_62_59 = p_62_61 & p_60_59;
 assign g_62_59 = g_62_61 | (p_62_61 & g_60_59);
 assign p_62_60 = p_62_61 & p_60_60;
 assign g_62_60 = g_62_61 | (p_62_61 & g_60_60);
 assign p_62_61 = p_62_62 & p_61_61;
 assign g_62_61 = g_62_62 | (p_62_62 & g_61_61);
 assign sum[62] = p_62_62^ g_61_0;
 assign cout = g_62_0;
endmodule
