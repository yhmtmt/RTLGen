module MG_CPA(
  input [31:0] a,
  input [31:0] b,
  output [31:0] sum,
  output cout
);

  wire p_0_0;
  wire g_0_0;
 assign p_0_0 = a[0] ^ b[0];
 assign g_0_0 = a[0] & b[0];
  wire p_1_1;
  wire g_1_1;
 assign p_1_1 = a[1] ^ b[1];
 assign g_1_1 = a[1] & b[1];
  wire p_1_0;
  wire g_1_0;
  wire p_2_2;
  wire g_2_2;
 assign p_2_2 = a[2] ^ b[2];
 assign g_2_2 = a[2] & b[2];
  wire p_2_0;
  wire g_2_0;
  wire p_3_3;
  wire g_3_3;
 assign p_3_3 = a[3] ^ b[3];
 assign g_3_3 = a[3] & b[3];
  wire p_3_0;
  wire g_3_0;
  wire p_3_2;
  wire g_3_2;
  wire p_4_4;
  wire g_4_4;
 assign p_4_4 = a[4] ^ b[4];
 assign g_4_4 = a[4] & b[4];
  wire p_4_0;
  wire g_4_0;
  wire p_5_5;
  wire g_5_5;
 assign p_5_5 = a[5] ^ b[5];
 assign g_5_5 = a[5] & b[5];
  wire p_5_0;
  wire g_5_0;
  wire p_5_4;
  wire g_5_4;
  wire p_6_6;
  wire g_6_6;
 assign p_6_6 = a[6] ^ b[6];
 assign g_6_6 = a[6] & b[6];
  wire p_6_0;
  wire g_6_0;
  wire p_7_7;
  wire g_7_7;
 assign p_7_7 = a[7] ^ b[7];
 assign g_7_7 = a[7] & b[7];
  wire p_7_0;
  wire g_7_0;
  wire p_7_4;
  wire g_7_4;
  wire p_7_6;
  wire g_7_6;
  wire p_8_8;
  wire g_8_8;
 assign p_8_8 = a[8] ^ b[8];
 assign g_8_8 = a[8] & b[8];
  wire p_8_0;
  wire g_8_0;
  wire p_9_9;
  wire g_9_9;
 assign p_9_9 = a[9] ^ b[9];
 assign g_9_9 = a[9] & b[9];
  wire p_9_0;
  wire g_9_0;
  wire p_9_8;
  wire g_9_8;
  wire p_10_10;
  wire g_10_10;
 assign p_10_10 = a[10] ^ b[10];
 assign g_10_10 = a[10] & b[10];
  wire p_10_0;
  wire g_10_0;
  wire p_11_11;
  wire g_11_11;
 assign p_11_11 = a[11] ^ b[11];
 assign g_11_11 = a[11] & b[11];
  wire p_11_0;
  wire g_11_0;
  wire p_11_8;
  wire g_11_8;
  wire p_11_10;
  wire g_11_10;
  wire p_12_12;
  wire g_12_12;
 assign p_12_12 = a[12] ^ b[12];
 assign g_12_12 = a[12] & b[12];
  wire p_12_0;
  wire g_12_0;
  wire p_13_13;
  wire g_13_13;
 assign p_13_13 = a[13] ^ b[13];
 assign g_13_13 = a[13] & b[13];
  wire p_13_0;
  wire g_13_0;
  wire p_13_12;
  wire g_13_12;
  wire p_14_14;
  wire g_14_14;
 assign p_14_14 = a[14] ^ b[14];
 assign g_14_14 = a[14] & b[14];
  wire p_14_0;
  wire g_14_0;
  wire p_15_15;
  wire g_15_15;
 assign p_15_15 = a[15] ^ b[15];
 assign g_15_15 = a[15] & b[15];
  wire p_15_0;
  wire g_15_0;
  wire p_15_8;
  wire g_15_8;
  wire p_15_12;
  wire g_15_12;
  wire p_15_14;
  wire g_15_14;
  wire p_16_16;
  wire g_16_16;
 assign p_16_16 = a[16] ^ b[16];
 assign g_16_16 = a[16] & b[16];
  wire p_16_0;
  wire g_16_0;
  wire p_17_17;
  wire g_17_17;
 assign p_17_17 = a[17] ^ b[17];
 assign g_17_17 = a[17] & b[17];
  wire p_17_0;
  wire g_17_0;
  wire p_17_16;
  wire g_17_16;
  wire p_18_18;
  wire g_18_18;
 assign p_18_18 = a[18] ^ b[18];
 assign g_18_18 = a[18] & b[18];
  wire p_18_0;
  wire g_18_0;
  wire p_19_19;
  wire g_19_19;
 assign p_19_19 = a[19] ^ b[19];
 assign g_19_19 = a[19] & b[19];
  wire p_19_0;
  wire g_19_0;
  wire p_19_16;
  wire g_19_16;
  wire p_19_18;
  wire g_19_18;
  wire p_20_20;
  wire g_20_20;
 assign p_20_20 = a[20] ^ b[20];
 assign g_20_20 = a[20] & b[20];
  wire p_20_0;
  wire g_20_0;
  wire p_21_21;
  wire g_21_21;
 assign p_21_21 = a[21] ^ b[21];
 assign g_21_21 = a[21] & b[21];
  wire p_21_0;
  wire g_21_0;
  wire p_21_20;
  wire g_21_20;
  wire p_22_22;
  wire g_22_22;
 assign p_22_22 = a[22] ^ b[22];
 assign g_22_22 = a[22] & b[22];
  wire p_22_0;
  wire g_22_0;
  wire p_23_23;
  wire g_23_23;
 assign p_23_23 = a[23] ^ b[23];
 assign g_23_23 = a[23] & b[23];
  wire p_23_0;
  wire g_23_0;
  wire p_23_16;
  wire g_23_16;
  wire p_23_20;
  wire g_23_20;
  wire p_23_22;
  wire g_23_22;
  wire p_24_24;
  wire g_24_24;
 assign p_24_24 = a[24] ^ b[24];
 assign g_24_24 = a[24] & b[24];
  wire p_24_0;
  wire g_24_0;
  wire p_25_25;
  wire g_25_25;
 assign p_25_25 = a[25] ^ b[25];
 assign g_25_25 = a[25] & b[25];
  wire p_25_0;
  wire g_25_0;
  wire p_25_24;
  wire g_25_24;
  wire p_26_26;
  wire g_26_26;
 assign p_26_26 = a[26] ^ b[26];
 assign g_26_26 = a[26] & b[26];
  wire p_26_0;
  wire g_26_0;
  wire p_27_27;
  wire g_27_27;
 assign p_27_27 = a[27] ^ b[27];
 assign g_27_27 = a[27] & b[27];
  wire p_27_0;
  wire g_27_0;
  wire p_27_24;
  wire g_27_24;
  wire p_27_26;
  wire g_27_26;
  wire p_28_28;
  wire g_28_28;
 assign p_28_28 = a[28] ^ b[28];
 assign g_28_28 = a[28] & b[28];
  wire p_28_0;
  wire g_28_0;
  wire p_29_29;
  wire g_29_29;
 assign p_29_29 = a[29] ^ b[29];
 assign g_29_29 = a[29] & b[29];
  wire p_29_0;
  wire g_29_0;
  wire p_29_28;
  wire g_29_28;
  wire p_30_30;
  wire g_30_30;
 assign p_30_30 = a[30] ^ b[30];
 assign g_30_30 = a[30] & b[30];
  wire p_30_0;
  wire g_30_0;
  wire p_31_31;
  wire g_31_31;
 assign p_31_31 = a[31] ^ b[31];
 assign g_31_31 = a[31] & b[31];
  wire p_31_0;
  wire g_31_0;
  wire p_31_16;
  wire g_31_16;
  wire p_31_24;
  wire g_31_24;
  wire p_31_28;
  wire g_31_28;
  wire p_31_30;
  wire g_31_30;
 assign sum[0] = p_0_0;
 assign p_1_0 = p_1_1 & p_0_0;
 assign g_1_0 = g_1_1 | (p_1_1 & g_0_0);
 assign sum[1] = p_1_1^ g_0_0;
 assign p_2_0 = p_2_2 & p_1_0;
 assign g_2_0 = g_2_2 | (p_2_2 & g_1_0);
 assign sum[2] = p_2_2^ g_1_0;
 assign p_3_0 = p_3_2 & p_1_0;
 assign g_3_0 = g_3_2 | (p_3_2 & g_1_0);
 assign p_3_2 = p_3_3 & p_2_2;
 assign g_3_2 = g_3_3 | (p_3_3 & g_2_2);
 assign sum[3] = p_3_3^ g_2_0;
 assign p_4_0 = p_4_4 & p_3_0;
 assign g_4_0 = g_4_4 | (p_4_4 & g_3_0);
 assign sum[4] = p_4_4^ g_3_0;
 assign p_5_0 = p_5_5 & p_4_0;
 assign g_5_0 = g_5_5 | (p_5_5 & g_4_0);
 assign p_5_4 = p_5_5 & p_4_4;
 assign g_5_4 = g_5_5 | (p_5_5 & g_4_4);
 assign sum[5] = p_5_5^ g_4_0;
 assign p_6_0 = p_6_6 & p_5_0;
 assign g_6_0 = g_6_6 | (p_6_6 & g_5_0);
 assign sum[6] = p_6_6^ g_5_0;
 assign p_7_0 = p_7_4 & p_3_0;
 assign g_7_0 = g_7_4 | (p_7_4 & g_3_0);
 assign p_7_4 = p_7_6 & p_5_4;
 assign g_7_4 = g_7_6 | (p_7_6 & g_5_4);
 assign p_7_6 = p_7_7 & p_6_6;
 assign g_7_6 = g_7_7 | (p_7_7 & g_6_6);
 assign sum[7] = p_7_7^ g_6_0;
 assign p_8_0 = p_8_8 & p_7_0;
 assign g_8_0 = g_8_8 | (p_8_8 & g_7_0);
 assign sum[8] = p_8_8^ g_7_0;
 assign p_9_0 = p_9_9 & p_8_0;
 assign g_9_0 = g_9_9 | (p_9_9 & g_8_0);
 assign p_9_8 = p_9_9 & p_8_8;
 assign g_9_8 = g_9_9 | (p_9_9 & g_8_8);
 assign sum[9] = p_9_9^ g_8_0;
 assign p_10_0 = p_10_10 & p_9_0;
 assign g_10_0 = g_10_10 | (p_10_10 & g_9_0);
 assign sum[10] = p_10_10^ g_9_0;
 assign p_11_0 = p_11_11 & p_10_0;
 assign g_11_0 = g_11_11 | (p_11_11 & g_10_0);
 assign p_11_8 = p_11_10 & p_9_8;
 assign g_11_8 = g_11_10 | (p_11_10 & g_9_8);
 assign p_11_10 = p_11_11 & p_10_10;
 assign g_11_10 = g_11_11 | (p_11_11 & g_10_10);
 assign sum[11] = p_11_11^ g_10_0;
 assign p_12_0 = p_12_12 & p_11_0;
 assign g_12_0 = g_12_12 | (p_12_12 & g_11_0);
 assign sum[12] = p_12_12^ g_11_0;
 assign p_13_0 = p_13_13 & p_12_0;
 assign g_13_0 = g_13_13 | (p_13_13 & g_12_0);
 assign p_13_12 = p_13_13 & p_12_12;
 assign g_13_12 = g_13_13 | (p_13_13 & g_12_12);
 assign sum[13] = p_13_13^ g_12_0;
 assign p_14_0 = p_14_14 & p_13_0;
 assign g_14_0 = g_14_14 | (p_14_14 & g_13_0);
 assign sum[14] = p_14_14^ g_13_0;
 assign p_15_0 = p_15_8 & p_7_0;
 assign g_15_0 = g_15_8 | (p_15_8 & g_7_0);
 assign p_15_8 = p_15_12 & p_11_8;
 assign g_15_8 = g_15_12 | (p_15_12 & g_11_8);
 assign p_15_12 = p_15_14 & p_13_12;
 assign g_15_12 = g_15_14 | (p_15_14 & g_13_12);
 assign p_15_14 = p_15_15 & p_14_14;
 assign g_15_14 = g_15_15 | (p_15_15 & g_14_14);
 assign sum[15] = p_15_15^ g_14_0;
 assign p_16_0 = p_16_16 & p_15_0;
 assign g_16_0 = g_16_16 | (p_16_16 & g_15_0);
 assign sum[16] = p_16_16^ g_15_0;
 assign p_17_0 = p_17_17 & p_16_0;
 assign g_17_0 = g_17_17 | (p_17_17 & g_16_0);
 assign p_17_16 = p_17_17 & p_16_16;
 assign g_17_16 = g_17_17 | (p_17_17 & g_16_16);
 assign sum[17] = p_17_17^ g_16_0;
 assign p_18_0 = p_18_18 & p_17_0;
 assign g_18_0 = g_18_18 | (p_18_18 & g_17_0);
 assign sum[18] = p_18_18^ g_17_0;
 assign p_19_0 = p_19_19 & p_18_0;
 assign g_19_0 = g_19_19 | (p_19_19 & g_18_0);
 assign p_19_16 = p_19_18 & p_17_16;
 assign g_19_16 = g_19_18 | (p_19_18 & g_17_16);
 assign p_19_18 = p_19_19 & p_18_18;
 assign g_19_18 = g_19_19 | (p_19_19 & g_18_18);
 assign sum[19] = p_19_19^ g_18_0;
 assign p_20_0 = p_20_20 & p_19_0;
 assign g_20_0 = g_20_20 | (p_20_20 & g_19_0);
 assign sum[20] = p_20_20^ g_19_0;
 assign p_21_0 = p_21_21 & p_20_0;
 assign g_21_0 = g_21_21 | (p_21_21 & g_20_0);
 assign p_21_20 = p_21_21 & p_20_20;
 assign g_21_20 = g_21_21 | (p_21_21 & g_20_20);
 assign sum[21] = p_21_21^ g_20_0;
 assign p_22_0 = p_22_22 & p_21_0;
 assign g_22_0 = g_22_22 | (p_22_22 & g_21_0);
 assign sum[22] = p_22_22^ g_21_0;
 assign p_23_0 = p_23_23 & p_22_0;
 assign g_23_0 = g_23_23 | (p_23_23 & g_22_0);
 assign p_23_16 = p_23_20 & p_19_16;
 assign g_23_16 = g_23_20 | (p_23_20 & g_19_16);
 assign p_23_20 = p_23_22 & p_21_20;
 assign g_23_20 = g_23_22 | (p_23_22 & g_21_20);
 assign p_23_22 = p_23_23 & p_22_22;
 assign g_23_22 = g_23_23 | (p_23_23 & g_22_22);
 assign sum[23] = p_23_23^ g_22_0;
 assign p_24_0 = p_24_24 & p_23_0;
 assign g_24_0 = g_24_24 | (p_24_24 & g_23_0);
 assign sum[24] = p_24_24^ g_23_0;
 assign p_25_0 = p_25_25 & p_24_0;
 assign g_25_0 = g_25_25 | (p_25_25 & g_24_0);
 assign p_25_24 = p_25_25 & p_24_24;
 assign g_25_24 = g_25_25 | (p_25_25 & g_24_24);
 assign sum[25] = p_25_25^ g_24_0;
 assign p_26_0 = p_26_26 & p_25_0;
 assign g_26_0 = g_26_26 | (p_26_26 & g_25_0);
 assign sum[26] = p_26_26^ g_25_0;
 assign p_27_0 = p_27_27 & p_26_0;
 assign g_27_0 = g_27_27 | (p_27_27 & g_26_0);
 assign p_27_24 = p_27_26 & p_25_24;
 assign g_27_24 = g_27_26 | (p_27_26 & g_25_24);
 assign p_27_26 = p_27_27 & p_26_26;
 assign g_27_26 = g_27_27 | (p_27_27 & g_26_26);
 assign sum[27] = p_27_27^ g_26_0;
 assign p_28_0 = p_28_28 & p_27_0;
 assign g_28_0 = g_28_28 | (p_28_28 & g_27_0);
 assign sum[28] = p_28_28^ g_27_0;
 assign p_29_0 = p_29_29 & p_28_0;
 assign g_29_0 = g_29_29 | (p_29_29 & g_28_0);
 assign p_29_28 = p_29_29 & p_28_28;
 assign g_29_28 = g_29_29 | (p_29_29 & g_28_28);
 assign sum[29] = p_29_29^ g_28_0;
 assign p_30_0 = p_30_30 & p_29_0;
 assign g_30_0 = g_30_30 | (p_30_30 & g_29_0);
 assign sum[30] = p_30_30^ g_29_0;
 assign p_31_0 = p_31_31 & p_30_0;
 assign g_31_0 = g_31_31 | (p_31_31 & g_30_0);
 assign p_31_16 = p_31_24 & p_23_16;
 assign g_31_16 = g_31_24 | (p_31_24 & g_23_16);
 assign p_31_24 = p_31_28 & p_27_24;
 assign g_31_24 = g_31_28 | (p_31_28 & g_27_24);
 assign p_31_28 = p_31_30 & p_29_28;
 assign g_31_28 = g_31_30 | (p_31_30 & g_29_28);
 assign p_31_30 = p_31_31 & p_30_30;
 assign g_31_30 = g_31_31 | (p_31_31 & g_30_30);
 assign sum[31] = p_31_31^ g_30_0;
 assign cout = g_31_0;
endmodule
