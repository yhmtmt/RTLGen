module MG_FA(
  input a,
  input b,
  input cin,
  output sum,
  output cout
);

  assign sum = (a ^ b) ^ cin;
  assign cout = (a & b) | (b & cin) | (a & cin);
endmodule
module MG_HA(
  input a,
  input b,
  output sum,
  output cout
);

  assign sum = a ^ b;
  assign cout = a & b;
endmodule
module mult32u_normal_sklansky(
  input [31:0] multiplicand,
  input [31:0] multiplier,
  output [63:0] product
);

  wire pp_0_0;
  wire pp_0_1;
  wire pp_0_10;
  wire pp_0_11;
  wire pp_0_12;
  wire pp_0_13;
  wire pp_0_14;
  wire pp_0_15;
  wire pp_0_16;
  wire pp_0_17;
  wire pp_0_18;
  wire pp_0_19;
  wire pp_0_2;
  wire pp_0_20;
  wire pp_0_21;
  wire pp_0_22;
  wire pp_0_23;
  wire pp_0_24;
  wire pp_0_25;
  wire pp_0_26;
  wire pp_0_27;
  wire pp_0_28;
  wire pp_0_29;
  wire pp_0_3;
  wire pp_0_30;
  wire pp_0_31;
  wire pp_0_4;
  wire pp_0_5;
  wire pp_0_6;
  wire pp_0_7;
  wire pp_0_8;
  wire pp_0_9;
  wire pp_10_10;
  wire pp_10_11;
  wire pp_10_12;
  wire pp_10_13;
  wire pp_10_14;
  wire pp_10_15;
  wire pp_10_16;
  wire pp_10_17;
  wire pp_10_18;
  wire pp_10_19;
  wire pp_10_20;
  wire pp_10_21;
  wire pp_10_22;
  wire pp_10_23;
  wire pp_10_24;
  wire pp_10_25;
  wire pp_10_26;
  wire pp_10_27;
  wire pp_10_28;
  wire pp_10_29;
  wire pp_10_30;
  wire pp_10_31;
  wire pp_10_32;
  wire pp_10_33;
  wire pp_10_34;
  wire pp_10_35;
  wire pp_10_36;
  wire pp_10_37;
  wire pp_10_38;
  wire pp_10_39;
  wire pp_10_40;
  wire pp_10_41;
  wire pp_11_11;
  wire pp_11_12;
  wire pp_11_13;
  wire pp_11_14;
  wire pp_11_15;
  wire pp_11_16;
  wire pp_11_17;
  wire pp_11_18;
  wire pp_11_19;
  wire pp_11_20;
  wire pp_11_21;
  wire pp_11_22;
  wire pp_11_23;
  wire pp_11_24;
  wire pp_11_25;
  wire pp_11_26;
  wire pp_11_27;
  wire pp_11_28;
  wire pp_11_29;
  wire pp_11_30;
  wire pp_11_31;
  wire pp_11_32;
  wire pp_11_33;
  wire pp_11_34;
  wire pp_11_35;
  wire pp_11_36;
  wire pp_11_37;
  wire pp_11_38;
  wire pp_11_39;
  wire pp_11_40;
  wire pp_11_41;
  wire pp_11_42;
  wire pp_12_12;
  wire pp_12_13;
  wire pp_12_14;
  wire pp_12_15;
  wire pp_12_16;
  wire pp_12_17;
  wire pp_12_18;
  wire pp_12_19;
  wire pp_12_20;
  wire pp_12_21;
  wire pp_12_22;
  wire pp_12_23;
  wire pp_12_24;
  wire pp_12_25;
  wire pp_12_26;
  wire pp_12_27;
  wire pp_12_28;
  wire pp_12_29;
  wire pp_12_30;
  wire pp_12_31;
  wire pp_12_32;
  wire pp_12_33;
  wire pp_12_34;
  wire pp_12_35;
  wire pp_12_36;
  wire pp_12_37;
  wire pp_12_38;
  wire pp_12_39;
  wire pp_12_40;
  wire pp_12_41;
  wire pp_12_42;
  wire pp_12_43;
  wire pp_13_13;
  wire pp_13_14;
  wire pp_13_15;
  wire pp_13_16;
  wire pp_13_17;
  wire pp_13_18;
  wire pp_13_19;
  wire pp_13_20;
  wire pp_13_21;
  wire pp_13_22;
  wire pp_13_23;
  wire pp_13_24;
  wire pp_13_25;
  wire pp_13_26;
  wire pp_13_27;
  wire pp_13_28;
  wire pp_13_29;
  wire pp_13_30;
  wire pp_13_31;
  wire pp_13_32;
  wire pp_13_33;
  wire pp_13_34;
  wire pp_13_35;
  wire pp_13_36;
  wire pp_13_37;
  wire pp_13_38;
  wire pp_13_39;
  wire pp_13_40;
  wire pp_13_41;
  wire pp_13_42;
  wire pp_13_43;
  wire pp_13_44;
  wire pp_14_14;
  wire pp_14_15;
  wire pp_14_16;
  wire pp_14_17;
  wire pp_14_18;
  wire pp_14_19;
  wire pp_14_20;
  wire pp_14_21;
  wire pp_14_22;
  wire pp_14_23;
  wire pp_14_24;
  wire pp_14_25;
  wire pp_14_26;
  wire pp_14_27;
  wire pp_14_28;
  wire pp_14_29;
  wire pp_14_30;
  wire pp_14_31;
  wire pp_14_32;
  wire pp_14_33;
  wire pp_14_34;
  wire pp_14_35;
  wire pp_14_36;
  wire pp_14_37;
  wire pp_14_38;
  wire pp_14_39;
  wire pp_14_40;
  wire pp_14_41;
  wire pp_14_42;
  wire pp_14_43;
  wire pp_14_44;
  wire pp_14_45;
  wire pp_15_15;
  wire pp_15_16;
  wire pp_15_17;
  wire pp_15_18;
  wire pp_15_19;
  wire pp_15_20;
  wire pp_15_21;
  wire pp_15_22;
  wire pp_15_23;
  wire pp_15_24;
  wire pp_15_25;
  wire pp_15_26;
  wire pp_15_27;
  wire pp_15_28;
  wire pp_15_29;
  wire pp_15_30;
  wire pp_15_31;
  wire pp_15_32;
  wire pp_15_33;
  wire pp_15_34;
  wire pp_15_35;
  wire pp_15_36;
  wire pp_15_37;
  wire pp_15_38;
  wire pp_15_39;
  wire pp_15_40;
  wire pp_15_41;
  wire pp_15_42;
  wire pp_15_43;
  wire pp_15_44;
  wire pp_15_45;
  wire pp_15_46;
  wire pp_16_16;
  wire pp_16_17;
  wire pp_16_18;
  wire pp_16_19;
  wire pp_16_20;
  wire pp_16_21;
  wire pp_16_22;
  wire pp_16_23;
  wire pp_16_24;
  wire pp_16_25;
  wire pp_16_26;
  wire pp_16_27;
  wire pp_16_28;
  wire pp_16_29;
  wire pp_16_30;
  wire pp_16_31;
  wire pp_16_32;
  wire pp_16_33;
  wire pp_16_34;
  wire pp_16_35;
  wire pp_16_36;
  wire pp_16_37;
  wire pp_16_38;
  wire pp_16_39;
  wire pp_16_40;
  wire pp_16_41;
  wire pp_16_42;
  wire pp_16_43;
  wire pp_16_44;
  wire pp_16_45;
  wire pp_16_46;
  wire pp_16_47;
  wire pp_17_17;
  wire pp_17_18;
  wire pp_17_19;
  wire pp_17_20;
  wire pp_17_21;
  wire pp_17_22;
  wire pp_17_23;
  wire pp_17_24;
  wire pp_17_25;
  wire pp_17_26;
  wire pp_17_27;
  wire pp_17_28;
  wire pp_17_29;
  wire pp_17_30;
  wire pp_17_31;
  wire pp_17_32;
  wire pp_17_33;
  wire pp_17_34;
  wire pp_17_35;
  wire pp_17_36;
  wire pp_17_37;
  wire pp_17_38;
  wire pp_17_39;
  wire pp_17_40;
  wire pp_17_41;
  wire pp_17_42;
  wire pp_17_43;
  wire pp_17_44;
  wire pp_17_45;
  wire pp_17_46;
  wire pp_17_47;
  wire pp_17_48;
  wire pp_18_18;
  wire pp_18_19;
  wire pp_18_20;
  wire pp_18_21;
  wire pp_18_22;
  wire pp_18_23;
  wire pp_18_24;
  wire pp_18_25;
  wire pp_18_26;
  wire pp_18_27;
  wire pp_18_28;
  wire pp_18_29;
  wire pp_18_30;
  wire pp_18_31;
  wire pp_18_32;
  wire pp_18_33;
  wire pp_18_34;
  wire pp_18_35;
  wire pp_18_36;
  wire pp_18_37;
  wire pp_18_38;
  wire pp_18_39;
  wire pp_18_40;
  wire pp_18_41;
  wire pp_18_42;
  wire pp_18_43;
  wire pp_18_44;
  wire pp_18_45;
  wire pp_18_46;
  wire pp_18_47;
  wire pp_18_48;
  wire pp_18_49;
  wire pp_19_19;
  wire pp_19_20;
  wire pp_19_21;
  wire pp_19_22;
  wire pp_19_23;
  wire pp_19_24;
  wire pp_19_25;
  wire pp_19_26;
  wire pp_19_27;
  wire pp_19_28;
  wire pp_19_29;
  wire pp_19_30;
  wire pp_19_31;
  wire pp_19_32;
  wire pp_19_33;
  wire pp_19_34;
  wire pp_19_35;
  wire pp_19_36;
  wire pp_19_37;
  wire pp_19_38;
  wire pp_19_39;
  wire pp_19_40;
  wire pp_19_41;
  wire pp_19_42;
  wire pp_19_43;
  wire pp_19_44;
  wire pp_19_45;
  wire pp_19_46;
  wire pp_19_47;
  wire pp_19_48;
  wire pp_19_49;
  wire pp_19_50;
  wire pp_1_1;
  wire pp_1_10;
  wire pp_1_11;
  wire pp_1_12;
  wire pp_1_13;
  wire pp_1_14;
  wire pp_1_15;
  wire pp_1_16;
  wire pp_1_17;
  wire pp_1_18;
  wire pp_1_19;
  wire pp_1_2;
  wire pp_1_20;
  wire pp_1_21;
  wire pp_1_22;
  wire pp_1_23;
  wire pp_1_24;
  wire pp_1_25;
  wire pp_1_26;
  wire pp_1_27;
  wire pp_1_28;
  wire pp_1_29;
  wire pp_1_3;
  wire pp_1_30;
  wire pp_1_31;
  wire pp_1_32;
  wire pp_1_4;
  wire pp_1_5;
  wire pp_1_6;
  wire pp_1_7;
  wire pp_1_8;
  wire pp_1_9;
  wire pp_20_20;
  wire pp_20_21;
  wire pp_20_22;
  wire pp_20_23;
  wire pp_20_24;
  wire pp_20_25;
  wire pp_20_26;
  wire pp_20_27;
  wire pp_20_28;
  wire pp_20_29;
  wire pp_20_30;
  wire pp_20_31;
  wire pp_20_32;
  wire pp_20_33;
  wire pp_20_34;
  wire pp_20_35;
  wire pp_20_36;
  wire pp_20_37;
  wire pp_20_38;
  wire pp_20_39;
  wire pp_20_40;
  wire pp_20_41;
  wire pp_20_42;
  wire pp_20_43;
  wire pp_20_44;
  wire pp_20_45;
  wire pp_20_46;
  wire pp_20_47;
  wire pp_20_48;
  wire pp_20_49;
  wire pp_20_50;
  wire pp_20_51;
  wire pp_21_21;
  wire pp_21_22;
  wire pp_21_23;
  wire pp_21_24;
  wire pp_21_25;
  wire pp_21_26;
  wire pp_21_27;
  wire pp_21_28;
  wire pp_21_29;
  wire pp_21_30;
  wire pp_21_31;
  wire pp_21_32;
  wire pp_21_33;
  wire pp_21_34;
  wire pp_21_35;
  wire pp_21_36;
  wire pp_21_37;
  wire pp_21_38;
  wire pp_21_39;
  wire pp_21_40;
  wire pp_21_41;
  wire pp_21_42;
  wire pp_21_43;
  wire pp_21_44;
  wire pp_21_45;
  wire pp_21_46;
  wire pp_21_47;
  wire pp_21_48;
  wire pp_21_49;
  wire pp_21_50;
  wire pp_21_51;
  wire pp_21_52;
  wire pp_22_22;
  wire pp_22_23;
  wire pp_22_24;
  wire pp_22_25;
  wire pp_22_26;
  wire pp_22_27;
  wire pp_22_28;
  wire pp_22_29;
  wire pp_22_30;
  wire pp_22_31;
  wire pp_22_32;
  wire pp_22_33;
  wire pp_22_34;
  wire pp_22_35;
  wire pp_22_36;
  wire pp_22_37;
  wire pp_22_38;
  wire pp_22_39;
  wire pp_22_40;
  wire pp_22_41;
  wire pp_22_42;
  wire pp_22_43;
  wire pp_22_44;
  wire pp_22_45;
  wire pp_22_46;
  wire pp_22_47;
  wire pp_22_48;
  wire pp_22_49;
  wire pp_22_50;
  wire pp_22_51;
  wire pp_22_52;
  wire pp_22_53;
  wire pp_23_23;
  wire pp_23_24;
  wire pp_23_25;
  wire pp_23_26;
  wire pp_23_27;
  wire pp_23_28;
  wire pp_23_29;
  wire pp_23_30;
  wire pp_23_31;
  wire pp_23_32;
  wire pp_23_33;
  wire pp_23_34;
  wire pp_23_35;
  wire pp_23_36;
  wire pp_23_37;
  wire pp_23_38;
  wire pp_23_39;
  wire pp_23_40;
  wire pp_23_41;
  wire pp_23_42;
  wire pp_23_43;
  wire pp_23_44;
  wire pp_23_45;
  wire pp_23_46;
  wire pp_23_47;
  wire pp_23_48;
  wire pp_23_49;
  wire pp_23_50;
  wire pp_23_51;
  wire pp_23_52;
  wire pp_23_53;
  wire pp_23_54;
  wire pp_24_24;
  wire pp_24_25;
  wire pp_24_26;
  wire pp_24_27;
  wire pp_24_28;
  wire pp_24_29;
  wire pp_24_30;
  wire pp_24_31;
  wire pp_24_32;
  wire pp_24_33;
  wire pp_24_34;
  wire pp_24_35;
  wire pp_24_36;
  wire pp_24_37;
  wire pp_24_38;
  wire pp_24_39;
  wire pp_24_40;
  wire pp_24_41;
  wire pp_24_42;
  wire pp_24_43;
  wire pp_24_44;
  wire pp_24_45;
  wire pp_24_46;
  wire pp_24_47;
  wire pp_24_48;
  wire pp_24_49;
  wire pp_24_50;
  wire pp_24_51;
  wire pp_24_52;
  wire pp_24_53;
  wire pp_24_54;
  wire pp_24_55;
  wire pp_25_25;
  wire pp_25_26;
  wire pp_25_27;
  wire pp_25_28;
  wire pp_25_29;
  wire pp_25_30;
  wire pp_25_31;
  wire pp_25_32;
  wire pp_25_33;
  wire pp_25_34;
  wire pp_25_35;
  wire pp_25_36;
  wire pp_25_37;
  wire pp_25_38;
  wire pp_25_39;
  wire pp_25_40;
  wire pp_25_41;
  wire pp_25_42;
  wire pp_25_43;
  wire pp_25_44;
  wire pp_25_45;
  wire pp_25_46;
  wire pp_25_47;
  wire pp_25_48;
  wire pp_25_49;
  wire pp_25_50;
  wire pp_25_51;
  wire pp_25_52;
  wire pp_25_53;
  wire pp_25_54;
  wire pp_25_55;
  wire pp_25_56;
  wire pp_26_26;
  wire pp_26_27;
  wire pp_26_28;
  wire pp_26_29;
  wire pp_26_30;
  wire pp_26_31;
  wire pp_26_32;
  wire pp_26_33;
  wire pp_26_34;
  wire pp_26_35;
  wire pp_26_36;
  wire pp_26_37;
  wire pp_26_38;
  wire pp_26_39;
  wire pp_26_40;
  wire pp_26_41;
  wire pp_26_42;
  wire pp_26_43;
  wire pp_26_44;
  wire pp_26_45;
  wire pp_26_46;
  wire pp_26_47;
  wire pp_26_48;
  wire pp_26_49;
  wire pp_26_50;
  wire pp_26_51;
  wire pp_26_52;
  wire pp_26_53;
  wire pp_26_54;
  wire pp_26_55;
  wire pp_26_56;
  wire pp_26_57;
  wire pp_27_27;
  wire pp_27_28;
  wire pp_27_29;
  wire pp_27_30;
  wire pp_27_31;
  wire pp_27_32;
  wire pp_27_33;
  wire pp_27_34;
  wire pp_27_35;
  wire pp_27_36;
  wire pp_27_37;
  wire pp_27_38;
  wire pp_27_39;
  wire pp_27_40;
  wire pp_27_41;
  wire pp_27_42;
  wire pp_27_43;
  wire pp_27_44;
  wire pp_27_45;
  wire pp_27_46;
  wire pp_27_47;
  wire pp_27_48;
  wire pp_27_49;
  wire pp_27_50;
  wire pp_27_51;
  wire pp_27_52;
  wire pp_27_53;
  wire pp_27_54;
  wire pp_27_55;
  wire pp_27_56;
  wire pp_27_57;
  wire pp_27_58;
  wire pp_28_28;
  wire pp_28_29;
  wire pp_28_30;
  wire pp_28_31;
  wire pp_28_32;
  wire pp_28_33;
  wire pp_28_34;
  wire pp_28_35;
  wire pp_28_36;
  wire pp_28_37;
  wire pp_28_38;
  wire pp_28_39;
  wire pp_28_40;
  wire pp_28_41;
  wire pp_28_42;
  wire pp_28_43;
  wire pp_28_44;
  wire pp_28_45;
  wire pp_28_46;
  wire pp_28_47;
  wire pp_28_48;
  wire pp_28_49;
  wire pp_28_50;
  wire pp_28_51;
  wire pp_28_52;
  wire pp_28_53;
  wire pp_28_54;
  wire pp_28_55;
  wire pp_28_56;
  wire pp_28_57;
  wire pp_28_58;
  wire pp_28_59;
  wire pp_29_29;
  wire pp_29_30;
  wire pp_29_31;
  wire pp_29_32;
  wire pp_29_33;
  wire pp_29_34;
  wire pp_29_35;
  wire pp_29_36;
  wire pp_29_37;
  wire pp_29_38;
  wire pp_29_39;
  wire pp_29_40;
  wire pp_29_41;
  wire pp_29_42;
  wire pp_29_43;
  wire pp_29_44;
  wire pp_29_45;
  wire pp_29_46;
  wire pp_29_47;
  wire pp_29_48;
  wire pp_29_49;
  wire pp_29_50;
  wire pp_29_51;
  wire pp_29_52;
  wire pp_29_53;
  wire pp_29_54;
  wire pp_29_55;
  wire pp_29_56;
  wire pp_29_57;
  wire pp_29_58;
  wire pp_29_59;
  wire pp_29_60;
  wire pp_2_10;
  wire pp_2_11;
  wire pp_2_12;
  wire pp_2_13;
  wire pp_2_14;
  wire pp_2_15;
  wire pp_2_16;
  wire pp_2_17;
  wire pp_2_18;
  wire pp_2_19;
  wire pp_2_2;
  wire pp_2_20;
  wire pp_2_21;
  wire pp_2_22;
  wire pp_2_23;
  wire pp_2_24;
  wire pp_2_25;
  wire pp_2_26;
  wire pp_2_27;
  wire pp_2_28;
  wire pp_2_29;
  wire pp_2_3;
  wire pp_2_30;
  wire pp_2_31;
  wire pp_2_32;
  wire pp_2_33;
  wire pp_2_4;
  wire pp_2_5;
  wire pp_2_6;
  wire pp_2_7;
  wire pp_2_8;
  wire pp_2_9;
  wire pp_30_30;
  wire pp_30_31;
  wire pp_30_32;
  wire pp_30_33;
  wire pp_30_34;
  wire pp_30_35;
  wire pp_30_36;
  wire pp_30_37;
  wire pp_30_38;
  wire pp_30_39;
  wire pp_30_40;
  wire pp_30_41;
  wire pp_30_42;
  wire pp_30_43;
  wire pp_30_44;
  wire pp_30_45;
  wire pp_30_46;
  wire pp_30_47;
  wire pp_30_48;
  wire pp_30_49;
  wire pp_30_50;
  wire pp_30_51;
  wire pp_30_52;
  wire pp_30_53;
  wire pp_30_54;
  wire pp_30_55;
  wire pp_30_56;
  wire pp_30_57;
  wire pp_30_58;
  wire pp_30_59;
  wire pp_30_60;
  wire pp_30_61;
  wire pp_31_31;
  wire pp_31_32;
  wire pp_31_33;
  wire pp_31_34;
  wire pp_31_35;
  wire pp_31_36;
  wire pp_31_37;
  wire pp_31_38;
  wire pp_31_39;
  wire pp_31_40;
  wire pp_31_41;
  wire pp_31_42;
  wire pp_31_43;
  wire pp_31_44;
  wire pp_31_45;
  wire pp_31_46;
  wire pp_31_47;
  wire pp_31_48;
  wire pp_31_49;
  wire pp_31_50;
  wire pp_31_51;
  wire pp_31_52;
  wire pp_31_53;
  wire pp_31_54;
  wire pp_31_55;
  wire pp_31_56;
  wire pp_31_57;
  wire pp_31_58;
  wire pp_31_59;
  wire pp_31_60;
  wire pp_31_61;
  wire pp_31_62;
  wire pp_3_10;
  wire pp_3_11;
  wire pp_3_12;
  wire pp_3_13;
  wire pp_3_14;
  wire pp_3_15;
  wire pp_3_16;
  wire pp_3_17;
  wire pp_3_18;
  wire pp_3_19;
  wire pp_3_20;
  wire pp_3_21;
  wire pp_3_22;
  wire pp_3_23;
  wire pp_3_24;
  wire pp_3_25;
  wire pp_3_26;
  wire pp_3_27;
  wire pp_3_28;
  wire pp_3_29;
  wire pp_3_3;
  wire pp_3_30;
  wire pp_3_31;
  wire pp_3_32;
  wire pp_3_33;
  wire pp_3_34;
  wire pp_3_4;
  wire pp_3_5;
  wire pp_3_6;
  wire pp_3_7;
  wire pp_3_8;
  wire pp_3_9;
  wire pp_4_10;
  wire pp_4_11;
  wire pp_4_12;
  wire pp_4_13;
  wire pp_4_14;
  wire pp_4_15;
  wire pp_4_16;
  wire pp_4_17;
  wire pp_4_18;
  wire pp_4_19;
  wire pp_4_20;
  wire pp_4_21;
  wire pp_4_22;
  wire pp_4_23;
  wire pp_4_24;
  wire pp_4_25;
  wire pp_4_26;
  wire pp_4_27;
  wire pp_4_28;
  wire pp_4_29;
  wire pp_4_30;
  wire pp_4_31;
  wire pp_4_32;
  wire pp_4_33;
  wire pp_4_34;
  wire pp_4_35;
  wire pp_4_4;
  wire pp_4_5;
  wire pp_4_6;
  wire pp_4_7;
  wire pp_4_8;
  wire pp_4_9;
  wire pp_5_10;
  wire pp_5_11;
  wire pp_5_12;
  wire pp_5_13;
  wire pp_5_14;
  wire pp_5_15;
  wire pp_5_16;
  wire pp_5_17;
  wire pp_5_18;
  wire pp_5_19;
  wire pp_5_20;
  wire pp_5_21;
  wire pp_5_22;
  wire pp_5_23;
  wire pp_5_24;
  wire pp_5_25;
  wire pp_5_26;
  wire pp_5_27;
  wire pp_5_28;
  wire pp_5_29;
  wire pp_5_30;
  wire pp_5_31;
  wire pp_5_32;
  wire pp_5_33;
  wire pp_5_34;
  wire pp_5_35;
  wire pp_5_36;
  wire pp_5_5;
  wire pp_5_6;
  wire pp_5_7;
  wire pp_5_8;
  wire pp_5_9;
  wire pp_6_10;
  wire pp_6_11;
  wire pp_6_12;
  wire pp_6_13;
  wire pp_6_14;
  wire pp_6_15;
  wire pp_6_16;
  wire pp_6_17;
  wire pp_6_18;
  wire pp_6_19;
  wire pp_6_20;
  wire pp_6_21;
  wire pp_6_22;
  wire pp_6_23;
  wire pp_6_24;
  wire pp_6_25;
  wire pp_6_26;
  wire pp_6_27;
  wire pp_6_28;
  wire pp_6_29;
  wire pp_6_30;
  wire pp_6_31;
  wire pp_6_32;
  wire pp_6_33;
  wire pp_6_34;
  wire pp_6_35;
  wire pp_6_36;
  wire pp_6_37;
  wire pp_6_6;
  wire pp_6_7;
  wire pp_6_8;
  wire pp_6_9;
  wire pp_7_10;
  wire pp_7_11;
  wire pp_7_12;
  wire pp_7_13;
  wire pp_7_14;
  wire pp_7_15;
  wire pp_7_16;
  wire pp_7_17;
  wire pp_7_18;
  wire pp_7_19;
  wire pp_7_20;
  wire pp_7_21;
  wire pp_7_22;
  wire pp_7_23;
  wire pp_7_24;
  wire pp_7_25;
  wire pp_7_26;
  wire pp_7_27;
  wire pp_7_28;
  wire pp_7_29;
  wire pp_7_30;
  wire pp_7_31;
  wire pp_7_32;
  wire pp_7_33;
  wire pp_7_34;
  wire pp_7_35;
  wire pp_7_36;
  wire pp_7_37;
  wire pp_7_38;
  wire pp_7_7;
  wire pp_7_8;
  wire pp_7_9;
  wire pp_8_10;
  wire pp_8_11;
  wire pp_8_12;
  wire pp_8_13;
  wire pp_8_14;
  wire pp_8_15;
  wire pp_8_16;
  wire pp_8_17;
  wire pp_8_18;
  wire pp_8_19;
  wire pp_8_20;
  wire pp_8_21;
  wire pp_8_22;
  wire pp_8_23;
  wire pp_8_24;
  wire pp_8_25;
  wire pp_8_26;
  wire pp_8_27;
  wire pp_8_28;
  wire pp_8_29;
  wire pp_8_30;
  wire pp_8_31;
  wire pp_8_32;
  wire pp_8_33;
  wire pp_8_34;
  wire pp_8_35;
  wire pp_8_36;
  wire pp_8_37;
  wire pp_8_38;
  wire pp_8_39;
  wire pp_8_8;
  wire pp_8_9;
  wire pp_9_10;
  wire pp_9_11;
  wire pp_9_12;
  wire pp_9_13;
  wire pp_9_14;
  wire pp_9_15;
  wire pp_9_16;
  wire pp_9_17;
  wire pp_9_18;
  wire pp_9_19;
  wire pp_9_20;
  wire pp_9_21;
  wire pp_9_22;
  wire pp_9_23;
  wire pp_9_24;
  wire pp_9_25;
  wire pp_9_26;
  wire pp_9_27;
  wire pp_9_28;
  wire pp_9_29;
  wire pp_9_30;
  wire pp_9_31;
  wire pp_9_32;
  wire pp_9_33;
  wire pp_9_34;
  wire pp_9_35;
  wire pp_9_36;
  wire pp_9_37;
  wire pp_9_38;
  wire pp_9_39;
  wire pp_9_40;
  wire pp_9_9;
  assign pp_0_0 = multiplicand[0] & multiplier[0];
  assign pp_0_1 = multiplicand[1] & multiplier[0];
  assign pp_0_10 = multiplicand[10] & multiplier[0];
  assign pp_0_11 = multiplicand[11] & multiplier[0];
  assign pp_0_12 = multiplicand[12] & multiplier[0];
  assign pp_0_13 = multiplicand[13] & multiplier[0];
  assign pp_0_14 = multiplicand[14] & multiplier[0];
  assign pp_0_15 = multiplicand[15] & multiplier[0];
  assign pp_0_16 = multiplicand[16] & multiplier[0];
  assign pp_0_17 = multiplicand[17] & multiplier[0];
  assign pp_0_18 = multiplicand[18] & multiplier[0];
  assign pp_0_19 = multiplicand[19] & multiplier[0];
  assign pp_0_2 = multiplicand[2] & multiplier[0];
  assign pp_0_20 = multiplicand[20] & multiplier[0];
  assign pp_0_21 = multiplicand[21] & multiplier[0];
  assign pp_0_22 = multiplicand[22] & multiplier[0];
  assign pp_0_23 = multiplicand[23] & multiplier[0];
  assign pp_0_24 = multiplicand[24] & multiplier[0];
  assign pp_0_25 = multiplicand[25] & multiplier[0];
  assign pp_0_26 = multiplicand[26] & multiplier[0];
  assign pp_0_27 = multiplicand[27] & multiplier[0];
  assign pp_0_28 = multiplicand[28] & multiplier[0];
  assign pp_0_29 = multiplicand[29] & multiplier[0];
  assign pp_0_3 = multiplicand[3] & multiplier[0];
  assign pp_0_30 = multiplicand[30] & multiplier[0];
  assign pp_0_31 = multiplicand[31] & multiplier[0];
  assign pp_0_4 = multiplicand[4] & multiplier[0];
  assign pp_0_5 = multiplicand[5] & multiplier[0];
  assign pp_0_6 = multiplicand[6] & multiplier[0];
  assign pp_0_7 = multiplicand[7] & multiplier[0];
  assign pp_0_8 = multiplicand[8] & multiplier[0];
  assign pp_0_9 = multiplicand[9] & multiplier[0];
  assign pp_10_10 = multiplicand[0] & multiplier[10];
  assign pp_10_11 = multiplicand[1] & multiplier[10];
  assign pp_10_12 = multiplicand[2] & multiplier[10];
  assign pp_10_13 = multiplicand[3] & multiplier[10];
  assign pp_10_14 = multiplicand[4] & multiplier[10];
  assign pp_10_15 = multiplicand[5] & multiplier[10];
  assign pp_10_16 = multiplicand[6] & multiplier[10];
  assign pp_10_17 = multiplicand[7] & multiplier[10];
  assign pp_10_18 = multiplicand[8] & multiplier[10];
  assign pp_10_19 = multiplicand[9] & multiplier[10];
  assign pp_10_20 = multiplicand[10] & multiplier[10];
  assign pp_10_21 = multiplicand[11] & multiplier[10];
  assign pp_10_22 = multiplicand[12] & multiplier[10];
  assign pp_10_23 = multiplicand[13] & multiplier[10];
  assign pp_10_24 = multiplicand[14] & multiplier[10];
  assign pp_10_25 = multiplicand[15] & multiplier[10];
  assign pp_10_26 = multiplicand[16] & multiplier[10];
  assign pp_10_27 = multiplicand[17] & multiplier[10];
  assign pp_10_28 = multiplicand[18] & multiplier[10];
  assign pp_10_29 = multiplicand[19] & multiplier[10];
  assign pp_10_30 = multiplicand[20] & multiplier[10];
  assign pp_10_31 = multiplicand[21] & multiplier[10];
  assign pp_10_32 = multiplicand[22] & multiplier[10];
  assign pp_10_33 = multiplicand[23] & multiplier[10];
  assign pp_10_34 = multiplicand[24] & multiplier[10];
  assign pp_10_35 = multiplicand[25] & multiplier[10];
  assign pp_10_36 = multiplicand[26] & multiplier[10];
  assign pp_10_37 = multiplicand[27] & multiplier[10];
  assign pp_10_38 = multiplicand[28] & multiplier[10];
  assign pp_10_39 = multiplicand[29] & multiplier[10];
  assign pp_10_40 = multiplicand[30] & multiplier[10];
  assign pp_10_41 = multiplicand[31] & multiplier[10];
  assign pp_11_11 = multiplicand[0] & multiplier[11];
  assign pp_11_12 = multiplicand[1] & multiplier[11];
  assign pp_11_13 = multiplicand[2] & multiplier[11];
  assign pp_11_14 = multiplicand[3] & multiplier[11];
  assign pp_11_15 = multiplicand[4] & multiplier[11];
  assign pp_11_16 = multiplicand[5] & multiplier[11];
  assign pp_11_17 = multiplicand[6] & multiplier[11];
  assign pp_11_18 = multiplicand[7] & multiplier[11];
  assign pp_11_19 = multiplicand[8] & multiplier[11];
  assign pp_11_20 = multiplicand[9] & multiplier[11];
  assign pp_11_21 = multiplicand[10] & multiplier[11];
  assign pp_11_22 = multiplicand[11] & multiplier[11];
  assign pp_11_23 = multiplicand[12] & multiplier[11];
  assign pp_11_24 = multiplicand[13] & multiplier[11];
  assign pp_11_25 = multiplicand[14] & multiplier[11];
  assign pp_11_26 = multiplicand[15] & multiplier[11];
  assign pp_11_27 = multiplicand[16] & multiplier[11];
  assign pp_11_28 = multiplicand[17] & multiplier[11];
  assign pp_11_29 = multiplicand[18] & multiplier[11];
  assign pp_11_30 = multiplicand[19] & multiplier[11];
  assign pp_11_31 = multiplicand[20] & multiplier[11];
  assign pp_11_32 = multiplicand[21] & multiplier[11];
  assign pp_11_33 = multiplicand[22] & multiplier[11];
  assign pp_11_34 = multiplicand[23] & multiplier[11];
  assign pp_11_35 = multiplicand[24] & multiplier[11];
  assign pp_11_36 = multiplicand[25] & multiplier[11];
  assign pp_11_37 = multiplicand[26] & multiplier[11];
  assign pp_11_38 = multiplicand[27] & multiplier[11];
  assign pp_11_39 = multiplicand[28] & multiplier[11];
  assign pp_11_40 = multiplicand[29] & multiplier[11];
  assign pp_11_41 = multiplicand[30] & multiplier[11];
  assign pp_11_42 = multiplicand[31] & multiplier[11];
  assign pp_12_12 = multiplicand[0] & multiplier[12];
  assign pp_12_13 = multiplicand[1] & multiplier[12];
  assign pp_12_14 = multiplicand[2] & multiplier[12];
  assign pp_12_15 = multiplicand[3] & multiplier[12];
  assign pp_12_16 = multiplicand[4] & multiplier[12];
  assign pp_12_17 = multiplicand[5] & multiplier[12];
  assign pp_12_18 = multiplicand[6] & multiplier[12];
  assign pp_12_19 = multiplicand[7] & multiplier[12];
  assign pp_12_20 = multiplicand[8] & multiplier[12];
  assign pp_12_21 = multiplicand[9] & multiplier[12];
  assign pp_12_22 = multiplicand[10] & multiplier[12];
  assign pp_12_23 = multiplicand[11] & multiplier[12];
  assign pp_12_24 = multiplicand[12] & multiplier[12];
  assign pp_12_25 = multiplicand[13] & multiplier[12];
  assign pp_12_26 = multiplicand[14] & multiplier[12];
  assign pp_12_27 = multiplicand[15] & multiplier[12];
  assign pp_12_28 = multiplicand[16] & multiplier[12];
  assign pp_12_29 = multiplicand[17] & multiplier[12];
  assign pp_12_30 = multiplicand[18] & multiplier[12];
  assign pp_12_31 = multiplicand[19] & multiplier[12];
  assign pp_12_32 = multiplicand[20] & multiplier[12];
  assign pp_12_33 = multiplicand[21] & multiplier[12];
  assign pp_12_34 = multiplicand[22] & multiplier[12];
  assign pp_12_35 = multiplicand[23] & multiplier[12];
  assign pp_12_36 = multiplicand[24] & multiplier[12];
  assign pp_12_37 = multiplicand[25] & multiplier[12];
  assign pp_12_38 = multiplicand[26] & multiplier[12];
  assign pp_12_39 = multiplicand[27] & multiplier[12];
  assign pp_12_40 = multiplicand[28] & multiplier[12];
  assign pp_12_41 = multiplicand[29] & multiplier[12];
  assign pp_12_42 = multiplicand[30] & multiplier[12];
  assign pp_12_43 = multiplicand[31] & multiplier[12];
  assign pp_13_13 = multiplicand[0] & multiplier[13];
  assign pp_13_14 = multiplicand[1] & multiplier[13];
  assign pp_13_15 = multiplicand[2] & multiplier[13];
  assign pp_13_16 = multiplicand[3] & multiplier[13];
  assign pp_13_17 = multiplicand[4] & multiplier[13];
  assign pp_13_18 = multiplicand[5] & multiplier[13];
  assign pp_13_19 = multiplicand[6] & multiplier[13];
  assign pp_13_20 = multiplicand[7] & multiplier[13];
  assign pp_13_21 = multiplicand[8] & multiplier[13];
  assign pp_13_22 = multiplicand[9] & multiplier[13];
  assign pp_13_23 = multiplicand[10] & multiplier[13];
  assign pp_13_24 = multiplicand[11] & multiplier[13];
  assign pp_13_25 = multiplicand[12] & multiplier[13];
  assign pp_13_26 = multiplicand[13] & multiplier[13];
  assign pp_13_27 = multiplicand[14] & multiplier[13];
  assign pp_13_28 = multiplicand[15] & multiplier[13];
  assign pp_13_29 = multiplicand[16] & multiplier[13];
  assign pp_13_30 = multiplicand[17] & multiplier[13];
  assign pp_13_31 = multiplicand[18] & multiplier[13];
  assign pp_13_32 = multiplicand[19] & multiplier[13];
  assign pp_13_33 = multiplicand[20] & multiplier[13];
  assign pp_13_34 = multiplicand[21] & multiplier[13];
  assign pp_13_35 = multiplicand[22] & multiplier[13];
  assign pp_13_36 = multiplicand[23] & multiplier[13];
  assign pp_13_37 = multiplicand[24] & multiplier[13];
  assign pp_13_38 = multiplicand[25] & multiplier[13];
  assign pp_13_39 = multiplicand[26] & multiplier[13];
  assign pp_13_40 = multiplicand[27] & multiplier[13];
  assign pp_13_41 = multiplicand[28] & multiplier[13];
  assign pp_13_42 = multiplicand[29] & multiplier[13];
  assign pp_13_43 = multiplicand[30] & multiplier[13];
  assign pp_13_44 = multiplicand[31] & multiplier[13];
  assign pp_14_14 = multiplicand[0] & multiplier[14];
  assign pp_14_15 = multiplicand[1] & multiplier[14];
  assign pp_14_16 = multiplicand[2] & multiplier[14];
  assign pp_14_17 = multiplicand[3] & multiplier[14];
  assign pp_14_18 = multiplicand[4] & multiplier[14];
  assign pp_14_19 = multiplicand[5] & multiplier[14];
  assign pp_14_20 = multiplicand[6] & multiplier[14];
  assign pp_14_21 = multiplicand[7] & multiplier[14];
  assign pp_14_22 = multiplicand[8] & multiplier[14];
  assign pp_14_23 = multiplicand[9] & multiplier[14];
  assign pp_14_24 = multiplicand[10] & multiplier[14];
  assign pp_14_25 = multiplicand[11] & multiplier[14];
  assign pp_14_26 = multiplicand[12] & multiplier[14];
  assign pp_14_27 = multiplicand[13] & multiplier[14];
  assign pp_14_28 = multiplicand[14] & multiplier[14];
  assign pp_14_29 = multiplicand[15] & multiplier[14];
  assign pp_14_30 = multiplicand[16] & multiplier[14];
  assign pp_14_31 = multiplicand[17] & multiplier[14];
  assign pp_14_32 = multiplicand[18] & multiplier[14];
  assign pp_14_33 = multiplicand[19] & multiplier[14];
  assign pp_14_34 = multiplicand[20] & multiplier[14];
  assign pp_14_35 = multiplicand[21] & multiplier[14];
  assign pp_14_36 = multiplicand[22] & multiplier[14];
  assign pp_14_37 = multiplicand[23] & multiplier[14];
  assign pp_14_38 = multiplicand[24] & multiplier[14];
  assign pp_14_39 = multiplicand[25] & multiplier[14];
  assign pp_14_40 = multiplicand[26] & multiplier[14];
  assign pp_14_41 = multiplicand[27] & multiplier[14];
  assign pp_14_42 = multiplicand[28] & multiplier[14];
  assign pp_14_43 = multiplicand[29] & multiplier[14];
  assign pp_14_44 = multiplicand[30] & multiplier[14];
  assign pp_14_45 = multiplicand[31] & multiplier[14];
  assign pp_15_15 = multiplicand[0] & multiplier[15];
  assign pp_15_16 = multiplicand[1] & multiplier[15];
  assign pp_15_17 = multiplicand[2] & multiplier[15];
  assign pp_15_18 = multiplicand[3] & multiplier[15];
  assign pp_15_19 = multiplicand[4] & multiplier[15];
  assign pp_15_20 = multiplicand[5] & multiplier[15];
  assign pp_15_21 = multiplicand[6] & multiplier[15];
  assign pp_15_22 = multiplicand[7] & multiplier[15];
  assign pp_15_23 = multiplicand[8] & multiplier[15];
  assign pp_15_24 = multiplicand[9] & multiplier[15];
  assign pp_15_25 = multiplicand[10] & multiplier[15];
  assign pp_15_26 = multiplicand[11] & multiplier[15];
  assign pp_15_27 = multiplicand[12] & multiplier[15];
  assign pp_15_28 = multiplicand[13] & multiplier[15];
  assign pp_15_29 = multiplicand[14] & multiplier[15];
  assign pp_15_30 = multiplicand[15] & multiplier[15];
  assign pp_15_31 = multiplicand[16] & multiplier[15];
  assign pp_15_32 = multiplicand[17] & multiplier[15];
  assign pp_15_33 = multiplicand[18] & multiplier[15];
  assign pp_15_34 = multiplicand[19] & multiplier[15];
  assign pp_15_35 = multiplicand[20] & multiplier[15];
  assign pp_15_36 = multiplicand[21] & multiplier[15];
  assign pp_15_37 = multiplicand[22] & multiplier[15];
  assign pp_15_38 = multiplicand[23] & multiplier[15];
  assign pp_15_39 = multiplicand[24] & multiplier[15];
  assign pp_15_40 = multiplicand[25] & multiplier[15];
  assign pp_15_41 = multiplicand[26] & multiplier[15];
  assign pp_15_42 = multiplicand[27] & multiplier[15];
  assign pp_15_43 = multiplicand[28] & multiplier[15];
  assign pp_15_44 = multiplicand[29] & multiplier[15];
  assign pp_15_45 = multiplicand[30] & multiplier[15];
  assign pp_15_46 = multiplicand[31] & multiplier[15];
  assign pp_16_16 = multiplicand[0] & multiplier[16];
  assign pp_16_17 = multiplicand[1] & multiplier[16];
  assign pp_16_18 = multiplicand[2] & multiplier[16];
  assign pp_16_19 = multiplicand[3] & multiplier[16];
  assign pp_16_20 = multiplicand[4] & multiplier[16];
  assign pp_16_21 = multiplicand[5] & multiplier[16];
  assign pp_16_22 = multiplicand[6] & multiplier[16];
  assign pp_16_23 = multiplicand[7] & multiplier[16];
  assign pp_16_24 = multiplicand[8] & multiplier[16];
  assign pp_16_25 = multiplicand[9] & multiplier[16];
  assign pp_16_26 = multiplicand[10] & multiplier[16];
  assign pp_16_27 = multiplicand[11] & multiplier[16];
  assign pp_16_28 = multiplicand[12] & multiplier[16];
  assign pp_16_29 = multiplicand[13] & multiplier[16];
  assign pp_16_30 = multiplicand[14] & multiplier[16];
  assign pp_16_31 = multiplicand[15] & multiplier[16];
  assign pp_16_32 = multiplicand[16] & multiplier[16];
  assign pp_16_33 = multiplicand[17] & multiplier[16];
  assign pp_16_34 = multiplicand[18] & multiplier[16];
  assign pp_16_35 = multiplicand[19] & multiplier[16];
  assign pp_16_36 = multiplicand[20] & multiplier[16];
  assign pp_16_37 = multiplicand[21] & multiplier[16];
  assign pp_16_38 = multiplicand[22] & multiplier[16];
  assign pp_16_39 = multiplicand[23] & multiplier[16];
  assign pp_16_40 = multiplicand[24] & multiplier[16];
  assign pp_16_41 = multiplicand[25] & multiplier[16];
  assign pp_16_42 = multiplicand[26] & multiplier[16];
  assign pp_16_43 = multiplicand[27] & multiplier[16];
  assign pp_16_44 = multiplicand[28] & multiplier[16];
  assign pp_16_45 = multiplicand[29] & multiplier[16];
  assign pp_16_46 = multiplicand[30] & multiplier[16];
  assign pp_16_47 = multiplicand[31] & multiplier[16];
  assign pp_17_17 = multiplicand[0] & multiplier[17];
  assign pp_17_18 = multiplicand[1] & multiplier[17];
  assign pp_17_19 = multiplicand[2] & multiplier[17];
  assign pp_17_20 = multiplicand[3] & multiplier[17];
  assign pp_17_21 = multiplicand[4] & multiplier[17];
  assign pp_17_22 = multiplicand[5] & multiplier[17];
  assign pp_17_23 = multiplicand[6] & multiplier[17];
  assign pp_17_24 = multiplicand[7] & multiplier[17];
  assign pp_17_25 = multiplicand[8] & multiplier[17];
  assign pp_17_26 = multiplicand[9] & multiplier[17];
  assign pp_17_27 = multiplicand[10] & multiplier[17];
  assign pp_17_28 = multiplicand[11] & multiplier[17];
  assign pp_17_29 = multiplicand[12] & multiplier[17];
  assign pp_17_30 = multiplicand[13] & multiplier[17];
  assign pp_17_31 = multiplicand[14] & multiplier[17];
  assign pp_17_32 = multiplicand[15] & multiplier[17];
  assign pp_17_33 = multiplicand[16] & multiplier[17];
  assign pp_17_34 = multiplicand[17] & multiplier[17];
  assign pp_17_35 = multiplicand[18] & multiplier[17];
  assign pp_17_36 = multiplicand[19] & multiplier[17];
  assign pp_17_37 = multiplicand[20] & multiplier[17];
  assign pp_17_38 = multiplicand[21] & multiplier[17];
  assign pp_17_39 = multiplicand[22] & multiplier[17];
  assign pp_17_40 = multiplicand[23] & multiplier[17];
  assign pp_17_41 = multiplicand[24] & multiplier[17];
  assign pp_17_42 = multiplicand[25] & multiplier[17];
  assign pp_17_43 = multiplicand[26] & multiplier[17];
  assign pp_17_44 = multiplicand[27] & multiplier[17];
  assign pp_17_45 = multiplicand[28] & multiplier[17];
  assign pp_17_46 = multiplicand[29] & multiplier[17];
  assign pp_17_47 = multiplicand[30] & multiplier[17];
  assign pp_17_48 = multiplicand[31] & multiplier[17];
  assign pp_18_18 = multiplicand[0] & multiplier[18];
  assign pp_18_19 = multiplicand[1] & multiplier[18];
  assign pp_18_20 = multiplicand[2] & multiplier[18];
  assign pp_18_21 = multiplicand[3] & multiplier[18];
  assign pp_18_22 = multiplicand[4] & multiplier[18];
  assign pp_18_23 = multiplicand[5] & multiplier[18];
  assign pp_18_24 = multiplicand[6] & multiplier[18];
  assign pp_18_25 = multiplicand[7] & multiplier[18];
  assign pp_18_26 = multiplicand[8] & multiplier[18];
  assign pp_18_27 = multiplicand[9] & multiplier[18];
  assign pp_18_28 = multiplicand[10] & multiplier[18];
  assign pp_18_29 = multiplicand[11] & multiplier[18];
  assign pp_18_30 = multiplicand[12] & multiplier[18];
  assign pp_18_31 = multiplicand[13] & multiplier[18];
  assign pp_18_32 = multiplicand[14] & multiplier[18];
  assign pp_18_33 = multiplicand[15] & multiplier[18];
  assign pp_18_34 = multiplicand[16] & multiplier[18];
  assign pp_18_35 = multiplicand[17] & multiplier[18];
  assign pp_18_36 = multiplicand[18] & multiplier[18];
  assign pp_18_37 = multiplicand[19] & multiplier[18];
  assign pp_18_38 = multiplicand[20] & multiplier[18];
  assign pp_18_39 = multiplicand[21] & multiplier[18];
  assign pp_18_40 = multiplicand[22] & multiplier[18];
  assign pp_18_41 = multiplicand[23] & multiplier[18];
  assign pp_18_42 = multiplicand[24] & multiplier[18];
  assign pp_18_43 = multiplicand[25] & multiplier[18];
  assign pp_18_44 = multiplicand[26] & multiplier[18];
  assign pp_18_45 = multiplicand[27] & multiplier[18];
  assign pp_18_46 = multiplicand[28] & multiplier[18];
  assign pp_18_47 = multiplicand[29] & multiplier[18];
  assign pp_18_48 = multiplicand[30] & multiplier[18];
  assign pp_18_49 = multiplicand[31] & multiplier[18];
  assign pp_19_19 = multiplicand[0] & multiplier[19];
  assign pp_19_20 = multiplicand[1] & multiplier[19];
  assign pp_19_21 = multiplicand[2] & multiplier[19];
  assign pp_19_22 = multiplicand[3] & multiplier[19];
  assign pp_19_23 = multiplicand[4] & multiplier[19];
  assign pp_19_24 = multiplicand[5] & multiplier[19];
  assign pp_19_25 = multiplicand[6] & multiplier[19];
  assign pp_19_26 = multiplicand[7] & multiplier[19];
  assign pp_19_27 = multiplicand[8] & multiplier[19];
  assign pp_19_28 = multiplicand[9] & multiplier[19];
  assign pp_19_29 = multiplicand[10] & multiplier[19];
  assign pp_19_30 = multiplicand[11] & multiplier[19];
  assign pp_19_31 = multiplicand[12] & multiplier[19];
  assign pp_19_32 = multiplicand[13] & multiplier[19];
  assign pp_19_33 = multiplicand[14] & multiplier[19];
  assign pp_19_34 = multiplicand[15] & multiplier[19];
  assign pp_19_35 = multiplicand[16] & multiplier[19];
  assign pp_19_36 = multiplicand[17] & multiplier[19];
  assign pp_19_37 = multiplicand[18] & multiplier[19];
  assign pp_19_38 = multiplicand[19] & multiplier[19];
  assign pp_19_39 = multiplicand[20] & multiplier[19];
  assign pp_19_40 = multiplicand[21] & multiplier[19];
  assign pp_19_41 = multiplicand[22] & multiplier[19];
  assign pp_19_42 = multiplicand[23] & multiplier[19];
  assign pp_19_43 = multiplicand[24] & multiplier[19];
  assign pp_19_44 = multiplicand[25] & multiplier[19];
  assign pp_19_45 = multiplicand[26] & multiplier[19];
  assign pp_19_46 = multiplicand[27] & multiplier[19];
  assign pp_19_47 = multiplicand[28] & multiplier[19];
  assign pp_19_48 = multiplicand[29] & multiplier[19];
  assign pp_19_49 = multiplicand[30] & multiplier[19];
  assign pp_19_50 = multiplicand[31] & multiplier[19];
  assign pp_1_1 = multiplicand[0] & multiplier[1];
  assign pp_1_10 = multiplicand[9] & multiplier[1];
  assign pp_1_11 = multiplicand[10] & multiplier[1];
  assign pp_1_12 = multiplicand[11] & multiplier[1];
  assign pp_1_13 = multiplicand[12] & multiplier[1];
  assign pp_1_14 = multiplicand[13] & multiplier[1];
  assign pp_1_15 = multiplicand[14] & multiplier[1];
  assign pp_1_16 = multiplicand[15] & multiplier[1];
  assign pp_1_17 = multiplicand[16] & multiplier[1];
  assign pp_1_18 = multiplicand[17] & multiplier[1];
  assign pp_1_19 = multiplicand[18] & multiplier[1];
  assign pp_1_2 = multiplicand[1] & multiplier[1];
  assign pp_1_20 = multiplicand[19] & multiplier[1];
  assign pp_1_21 = multiplicand[20] & multiplier[1];
  assign pp_1_22 = multiplicand[21] & multiplier[1];
  assign pp_1_23 = multiplicand[22] & multiplier[1];
  assign pp_1_24 = multiplicand[23] & multiplier[1];
  assign pp_1_25 = multiplicand[24] & multiplier[1];
  assign pp_1_26 = multiplicand[25] & multiplier[1];
  assign pp_1_27 = multiplicand[26] & multiplier[1];
  assign pp_1_28 = multiplicand[27] & multiplier[1];
  assign pp_1_29 = multiplicand[28] & multiplier[1];
  assign pp_1_3 = multiplicand[2] & multiplier[1];
  assign pp_1_30 = multiplicand[29] & multiplier[1];
  assign pp_1_31 = multiplicand[30] & multiplier[1];
  assign pp_1_32 = multiplicand[31] & multiplier[1];
  assign pp_1_4 = multiplicand[3] & multiplier[1];
  assign pp_1_5 = multiplicand[4] & multiplier[1];
  assign pp_1_6 = multiplicand[5] & multiplier[1];
  assign pp_1_7 = multiplicand[6] & multiplier[1];
  assign pp_1_8 = multiplicand[7] & multiplier[1];
  assign pp_1_9 = multiplicand[8] & multiplier[1];
  assign pp_20_20 = multiplicand[0] & multiplier[20];
  assign pp_20_21 = multiplicand[1] & multiplier[20];
  assign pp_20_22 = multiplicand[2] & multiplier[20];
  assign pp_20_23 = multiplicand[3] & multiplier[20];
  assign pp_20_24 = multiplicand[4] & multiplier[20];
  assign pp_20_25 = multiplicand[5] & multiplier[20];
  assign pp_20_26 = multiplicand[6] & multiplier[20];
  assign pp_20_27 = multiplicand[7] & multiplier[20];
  assign pp_20_28 = multiplicand[8] & multiplier[20];
  assign pp_20_29 = multiplicand[9] & multiplier[20];
  assign pp_20_30 = multiplicand[10] & multiplier[20];
  assign pp_20_31 = multiplicand[11] & multiplier[20];
  assign pp_20_32 = multiplicand[12] & multiplier[20];
  assign pp_20_33 = multiplicand[13] & multiplier[20];
  assign pp_20_34 = multiplicand[14] & multiplier[20];
  assign pp_20_35 = multiplicand[15] & multiplier[20];
  assign pp_20_36 = multiplicand[16] & multiplier[20];
  assign pp_20_37 = multiplicand[17] & multiplier[20];
  assign pp_20_38 = multiplicand[18] & multiplier[20];
  assign pp_20_39 = multiplicand[19] & multiplier[20];
  assign pp_20_40 = multiplicand[20] & multiplier[20];
  assign pp_20_41 = multiplicand[21] & multiplier[20];
  assign pp_20_42 = multiplicand[22] & multiplier[20];
  assign pp_20_43 = multiplicand[23] & multiplier[20];
  assign pp_20_44 = multiplicand[24] & multiplier[20];
  assign pp_20_45 = multiplicand[25] & multiplier[20];
  assign pp_20_46 = multiplicand[26] & multiplier[20];
  assign pp_20_47 = multiplicand[27] & multiplier[20];
  assign pp_20_48 = multiplicand[28] & multiplier[20];
  assign pp_20_49 = multiplicand[29] & multiplier[20];
  assign pp_20_50 = multiplicand[30] & multiplier[20];
  assign pp_20_51 = multiplicand[31] & multiplier[20];
  assign pp_21_21 = multiplicand[0] & multiplier[21];
  assign pp_21_22 = multiplicand[1] & multiplier[21];
  assign pp_21_23 = multiplicand[2] & multiplier[21];
  assign pp_21_24 = multiplicand[3] & multiplier[21];
  assign pp_21_25 = multiplicand[4] & multiplier[21];
  assign pp_21_26 = multiplicand[5] & multiplier[21];
  assign pp_21_27 = multiplicand[6] & multiplier[21];
  assign pp_21_28 = multiplicand[7] & multiplier[21];
  assign pp_21_29 = multiplicand[8] & multiplier[21];
  assign pp_21_30 = multiplicand[9] & multiplier[21];
  assign pp_21_31 = multiplicand[10] & multiplier[21];
  assign pp_21_32 = multiplicand[11] & multiplier[21];
  assign pp_21_33 = multiplicand[12] & multiplier[21];
  assign pp_21_34 = multiplicand[13] & multiplier[21];
  assign pp_21_35 = multiplicand[14] & multiplier[21];
  assign pp_21_36 = multiplicand[15] & multiplier[21];
  assign pp_21_37 = multiplicand[16] & multiplier[21];
  assign pp_21_38 = multiplicand[17] & multiplier[21];
  assign pp_21_39 = multiplicand[18] & multiplier[21];
  assign pp_21_40 = multiplicand[19] & multiplier[21];
  assign pp_21_41 = multiplicand[20] & multiplier[21];
  assign pp_21_42 = multiplicand[21] & multiplier[21];
  assign pp_21_43 = multiplicand[22] & multiplier[21];
  assign pp_21_44 = multiplicand[23] & multiplier[21];
  assign pp_21_45 = multiplicand[24] & multiplier[21];
  assign pp_21_46 = multiplicand[25] & multiplier[21];
  assign pp_21_47 = multiplicand[26] & multiplier[21];
  assign pp_21_48 = multiplicand[27] & multiplier[21];
  assign pp_21_49 = multiplicand[28] & multiplier[21];
  assign pp_21_50 = multiplicand[29] & multiplier[21];
  assign pp_21_51 = multiplicand[30] & multiplier[21];
  assign pp_21_52 = multiplicand[31] & multiplier[21];
  assign pp_22_22 = multiplicand[0] & multiplier[22];
  assign pp_22_23 = multiplicand[1] & multiplier[22];
  assign pp_22_24 = multiplicand[2] & multiplier[22];
  assign pp_22_25 = multiplicand[3] & multiplier[22];
  assign pp_22_26 = multiplicand[4] & multiplier[22];
  assign pp_22_27 = multiplicand[5] & multiplier[22];
  assign pp_22_28 = multiplicand[6] & multiplier[22];
  assign pp_22_29 = multiplicand[7] & multiplier[22];
  assign pp_22_30 = multiplicand[8] & multiplier[22];
  assign pp_22_31 = multiplicand[9] & multiplier[22];
  assign pp_22_32 = multiplicand[10] & multiplier[22];
  assign pp_22_33 = multiplicand[11] & multiplier[22];
  assign pp_22_34 = multiplicand[12] & multiplier[22];
  assign pp_22_35 = multiplicand[13] & multiplier[22];
  assign pp_22_36 = multiplicand[14] & multiplier[22];
  assign pp_22_37 = multiplicand[15] & multiplier[22];
  assign pp_22_38 = multiplicand[16] & multiplier[22];
  assign pp_22_39 = multiplicand[17] & multiplier[22];
  assign pp_22_40 = multiplicand[18] & multiplier[22];
  assign pp_22_41 = multiplicand[19] & multiplier[22];
  assign pp_22_42 = multiplicand[20] & multiplier[22];
  assign pp_22_43 = multiplicand[21] & multiplier[22];
  assign pp_22_44 = multiplicand[22] & multiplier[22];
  assign pp_22_45 = multiplicand[23] & multiplier[22];
  assign pp_22_46 = multiplicand[24] & multiplier[22];
  assign pp_22_47 = multiplicand[25] & multiplier[22];
  assign pp_22_48 = multiplicand[26] & multiplier[22];
  assign pp_22_49 = multiplicand[27] & multiplier[22];
  assign pp_22_50 = multiplicand[28] & multiplier[22];
  assign pp_22_51 = multiplicand[29] & multiplier[22];
  assign pp_22_52 = multiplicand[30] & multiplier[22];
  assign pp_22_53 = multiplicand[31] & multiplier[22];
  assign pp_23_23 = multiplicand[0] & multiplier[23];
  assign pp_23_24 = multiplicand[1] & multiplier[23];
  assign pp_23_25 = multiplicand[2] & multiplier[23];
  assign pp_23_26 = multiplicand[3] & multiplier[23];
  assign pp_23_27 = multiplicand[4] & multiplier[23];
  assign pp_23_28 = multiplicand[5] & multiplier[23];
  assign pp_23_29 = multiplicand[6] & multiplier[23];
  assign pp_23_30 = multiplicand[7] & multiplier[23];
  assign pp_23_31 = multiplicand[8] & multiplier[23];
  assign pp_23_32 = multiplicand[9] & multiplier[23];
  assign pp_23_33 = multiplicand[10] & multiplier[23];
  assign pp_23_34 = multiplicand[11] & multiplier[23];
  assign pp_23_35 = multiplicand[12] & multiplier[23];
  assign pp_23_36 = multiplicand[13] & multiplier[23];
  assign pp_23_37 = multiplicand[14] & multiplier[23];
  assign pp_23_38 = multiplicand[15] & multiplier[23];
  assign pp_23_39 = multiplicand[16] & multiplier[23];
  assign pp_23_40 = multiplicand[17] & multiplier[23];
  assign pp_23_41 = multiplicand[18] & multiplier[23];
  assign pp_23_42 = multiplicand[19] & multiplier[23];
  assign pp_23_43 = multiplicand[20] & multiplier[23];
  assign pp_23_44 = multiplicand[21] & multiplier[23];
  assign pp_23_45 = multiplicand[22] & multiplier[23];
  assign pp_23_46 = multiplicand[23] & multiplier[23];
  assign pp_23_47 = multiplicand[24] & multiplier[23];
  assign pp_23_48 = multiplicand[25] & multiplier[23];
  assign pp_23_49 = multiplicand[26] & multiplier[23];
  assign pp_23_50 = multiplicand[27] & multiplier[23];
  assign pp_23_51 = multiplicand[28] & multiplier[23];
  assign pp_23_52 = multiplicand[29] & multiplier[23];
  assign pp_23_53 = multiplicand[30] & multiplier[23];
  assign pp_23_54 = multiplicand[31] & multiplier[23];
  assign pp_24_24 = multiplicand[0] & multiplier[24];
  assign pp_24_25 = multiplicand[1] & multiplier[24];
  assign pp_24_26 = multiplicand[2] & multiplier[24];
  assign pp_24_27 = multiplicand[3] & multiplier[24];
  assign pp_24_28 = multiplicand[4] & multiplier[24];
  assign pp_24_29 = multiplicand[5] & multiplier[24];
  assign pp_24_30 = multiplicand[6] & multiplier[24];
  assign pp_24_31 = multiplicand[7] & multiplier[24];
  assign pp_24_32 = multiplicand[8] & multiplier[24];
  assign pp_24_33 = multiplicand[9] & multiplier[24];
  assign pp_24_34 = multiplicand[10] & multiplier[24];
  assign pp_24_35 = multiplicand[11] & multiplier[24];
  assign pp_24_36 = multiplicand[12] & multiplier[24];
  assign pp_24_37 = multiplicand[13] & multiplier[24];
  assign pp_24_38 = multiplicand[14] & multiplier[24];
  assign pp_24_39 = multiplicand[15] & multiplier[24];
  assign pp_24_40 = multiplicand[16] & multiplier[24];
  assign pp_24_41 = multiplicand[17] & multiplier[24];
  assign pp_24_42 = multiplicand[18] & multiplier[24];
  assign pp_24_43 = multiplicand[19] & multiplier[24];
  assign pp_24_44 = multiplicand[20] & multiplier[24];
  assign pp_24_45 = multiplicand[21] & multiplier[24];
  assign pp_24_46 = multiplicand[22] & multiplier[24];
  assign pp_24_47 = multiplicand[23] & multiplier[24];
  assign pp_24_48 = multiplicand[24] & multiplier[24];
  assign pp_24_49 = multiplicand[25] & multiplier[24];
  assign pp_24_50 = multiplicand[26] & multiplier[24];
  assign pp_24_51 = multiplicand[27] & multiplier[24];
  assign pp_24_52 = multiplicand[28] & multiplier[24];
  assign pp_24_53 = multiplicand[29] & multiplier[24];
  assign pp_24_54 = multiplicand[30] & multiplier[24];
  assign pp_24_55 = multiplicand[31] & multiplier[24];
  assign pp_25_25 = multiplicand[0] & multiplier[25];
  assign pp_25_26 = multiplicand[1] & multiplier[25];
  assign pp_25_27 = multiplicand[2] & multiplier[25];
  assign pp_25_28 = multiplicand[3] & multiplier[25];
  assign pp_25_29 = multiplicand[4] & multiplier[25];
  assign pp_25_30 = multiplicand[5] & multiplier[25];
  assign pp_25_31 = multiplicand[6] & multiplier[25];
  assign pp_25_32 = multiplicand[7] & multiplier[25];
  assign pp_25_33 = multiplicand[8] & multiplier[25];
  assign pp_25_34 = multiplicand[9] & multiplier[25];
  assign pp_25_35 = multiplicand[10] & multiplier[25];
  assign pp_25_36 = multiplicand[11] & multiplier[25];
  assign pp_25_37 = multiplicand[12] & multiplier[25];
  assign pp_25_38 = multiplicand[13] & multiplier[25];
  assign pp_25_39 = multiplicand[14] & multiplier[25];
  assign pp_25_40 = multiplicand[15] & multiplier[25];
  assign pp_25_41 = multiplicand[16] & multiplier[25];
  assign pp_25_42 = multiplicand[17] & multiplier[25];
  assign pp_25_43 = multiplicand[18] & multiplier[25];
  assign pp_25_44 = multiplicand[19] & multiplier[25];
  assign pp_25_45 = multiplicand[20] & multiplier[25];
  assign pp_25_46 = multiplicand[21] & multiplier[25];
  assign pp_25_47 = multiplicand[22] & multiplier[25];
  assign pp_25_48 = multiplicand[23] & multiplier[25];
  assign pp_25_49 = multiplicand[24] & multiplier[25];
  assign pp_25_50 = multiplicand[25] & multiplier[25];
  assign pp_25_51 = multiplicand[26] & multiplier[25];
  assign pp_25_52 = multiplicand[27] & multiplier[25];
  assign pp_25_53 = multiplicand[28] & multiplier[25];
  assign pp_25_54 = multiplicand[29] & multiplier[25];
  assign pp_25_55 = multiplicand[30] & multiplier[25];
  assign pp_25_56 = multiplicand[31] & multiplier[25];
  assign pp_26_26 = multiplicand[0] & multiplier[26];
  assign pp_26_27 = multiplicand[1] & multiplier[26];
  assign pp_26_28 = multiplicand[2] & multiplier[26];
  assign pp_26_29 = multiplicand[3] & multiplier[26];
  assign pp_26_30 = multiplicand[4] & multiplier[26];
  assign pp_26_31 = multiplicand[5] & multiplier[26];
  assign pp_26_32 = multiplicand[6] & multiplier[26];
  assign pp_26_33 = multiplicand[7] & multiplier[26];
  assign pp_26_34 = multiplicand[8] & multiplier[26];
  assign pp_26_35 = multiplicand[9] & multiplier[26];
  assign pp_26_36 = multiplicand[10] & multiplier[26];
  assign pp_26_37 = multiplicand[11] & multiplier[26];
  assign pp_26_38 = multiplicand[12] & multiplier[26];
  assign pp_26_39 = multiplicand[13] & multiplier[26];
  assign pp_26_40 = multiplicand[14] & multiplier[26];
  assign pp_26_41 = multiplicand[15] & multiplier[26];
  assign pp_26_42 = multiplicand[16] & multiplier[26];
  assign pp_26_43 = multiplicand[17] & multiplier[26];
  assign pp_26_44 = multiplicand[18] & multiplier[26];
  assign pp_26_45 = multiplicand[19] & multiplier[26];
  assign pp_26_46 = multiplicand[20] & multiplier[26];
  assign pp_26_47 = multiplicand[21] & multiplier[26];
  assign pp_26_48 = multiplicand[22] & multiplier[26];
  assign pp_26_49 = multiplicand[23] & multiplier[26];
  assign pp_26_50 = multiplicand[24] & multiplier[26];
  assign pp_26_51 = multiplicand[25] & multiplier[26];
  assign pp_26_52 = multiplicand[26] & multiplier[26];
  assign pp_26_53 = multiplicand[27] & multiplier[26];
  assign pp_26_54 = multiplicand[28] & multiplier[26];
  assign pp_26_55 = multiplicand[29] & multiplier[26];
  assign pp_26_56 = multiplicand[30] & multiplier[26];
  assign pp_26_57 = multiplicand[31] & multiplier[26];
  assign pp_27_27 = multiplicand[0] & multiplier[27];
  assign pp_27_28 = multiplicand[1] & multiplier[27];
  assign pp_27_29 = multiplicand[2] & multiplier[27];
  assign pp_27_30 = multiplicand[3] & multiplier[27];
  assign pp_27_31 = multiplicand[4] & multiplier[27];
  assign pp_27_32 = multiplicand[5] & multiplier[27];
  assign pp_27_33 = multiplicand[6] & multiplier[27];
  assign pp_27_34 = multiplicand[7] & multiplier[27];
  assign pp_27_35 = multiplicand[8] & multiplier[27];
  assign pp_27_36 = multiplicand[9] & multiplier[27];
  assign pp_27_37 = multiplicand[10] & multiplier[27];
  assign pp_27_38 = multiplicand[11] & multiplier[27];
  assign pp_27_39 = multiplicand[12] & multiplier[27];
  assign pp_27_40 = multiplicand[13] & multiplier[27];
  assign pp_27_41 = multiplicand[14] & multiplier[27];
  assign pp_27_42 = multiplicand[15] & multiplier[27];
  assign pp_27_43 = multiplicand[16] & multiplier[27];
  assign pp_27_44 = multiplicand[17] & multiplier[27];
  assign pp_27_45 = multiplicand[18] & multiplier[27];
  assign pp_27_46 = multiplicand[19] & multiplier[27];
  assign pp_27_47 = multiplicand[20] & multiplier[27];
  assign pp_27_48 = multiplicand[21] & multiplier[27];
  assign pp_27_49 = multiplicand[22] & multiplier[27];
  assign pp_27_50 = multiplicand[23] & multiplier[27];
  assign pp_27_51 = multiplicand[24] & multiplier[27];
  assign pp_27_52 = multiplicand[25] & multiplier[27];
  assign pp_27_53 = multiplicand[26] & multiplier[27];
  assign pp_27_54 = multiplicand[27] & multiplier[27];
  assign pp_27_55 = multiplicand[28] & multiplier[27];
  assign pp_27_56 = multiplicand[29] & multiplier[27];
  assign pp_27_57 = multiplicand[30] & multiplier[27];
  assign pp_27_58 = multiplicand[31] & multiplier[27];
  assign pp_28_28 = multiplicand[0] & multiplier[28];
  assign pp_28_29 = multiplicand[1] & multiplier[28];
  assign pp_28_30 = multiplicand[2] & multiplier[28];
  assign pp_28_31 = multiplicand[3] & multiplier[28];
  assign pp_28_32 = multiplicand[4] & multiplier[28];
  assign pp_28_33 = multiplicand[5] & multiplier[28];
  assign pp_28_34 = multiplicand[6] & multiplier[28];
  assign pp_28_35 = multiplicand[7] & multiplier[28];
  assign pp_28_36 = multiplicand[8] & multiplier[28];
  assign pp_28_37 = multiplicand[9] & multiplier[28];
  assign pp_28_38 = multiplicand[10] & multiplier[28];
  assign pp_28_39 = multiplicand[11] & multiplier[28];
  assign pp_28_40 = multiplicand[12] & multiplier[28];
  assign pp_28_41 = multiplicand[13] & multiplier[28];
  assign pp_28_42 = multiplicand[14] & multiplier[28];
  assign pp_28_43 = multiplicand[15] & multiplier[28];
  assign pp_28_44 = multiplicand[16] & multiplier[28];
  assign pp_28_45 = multiplicand[17] & multiplier[28];
  assign pp_28_46 = multiplicand[18] & multiplier[28];
  assign pp_28_47 = multiplicand[19] & multiplier[28];
  assign pp_28_48 = multiplicand[20] & multiplier[28];
  assign pp_28_49 = multiplicand[21] & multiplier[28];
  assign pp_28_50 = multiplicand[22] & multiplier[28];
  assign pp_28_51 = multiplicand[23] & multiplier[28];
  assign pp_28_52 = multiplicand[24] & multiplier[28];
  assign pp_28_53 = multiplicand[25] & multiplier[28];
  assign pp_28_54 = multiplicand[26] & multiplier[28];
  assign pp_28_55 = multiplicand[27] & multiplier[28];
  assign pp_28_56 = multiplicand[28] & multiplier[28];
  assign pp_28_57 = multiplicand[29] & multiplier[28];
  assign pp_28_58 = multiplicand[30] & multiplier[28];
  assign pp_28_59 = multiplicand[31] & multiplier[28];
  assign pp_29_29 = multiplicand[0] & multiplier[29];
  assign pp_29_30 = multiplicand[1] & multiplier[29];
  assign pp_29_31 = multiplicand[2] & multiplier[29];
  assign pp_29_32 = multiplicand[3] & multiplier[29];
  assign pp_29_33 = multiplicand[4] & multiplier[29];
  assign pp_29_34 = multiplicand[5] & multiplier[29];
  assign pp_29_35 = multiplicand[6] & multiplier[29];
  assign pp_29_36 = multiplicand[7] & multiplier[29];
  assign pp_29_37 = multiplicand[8] & multiplier[29];
  assign pp_29_38 = multiplicand[9] & multiplier[29];
  assign pp_29_39 = multiplicand[10] & multiplier[29];
  assign pp_29_40 = multiplicand[11] & multiplier[29];
  assign pp_29_41 = multiplicand[12] & multiplier[29];
  assign pp_29_42 = multiplicand[13] & multiplier[29];
  assign pp_29_43 = multiplicand[14] & multiplier[29];
  assign pp_29_44 = multiplicand[15] & multiplier[29];
  assign pp_29_45 = multiplicand[16] & multiplier[29];
  assign pp_29_46 = multiplicand[17] & multiplier[29];
  assign pp_29_47 = multiplicand[18] & multiplier[29];
  assign pp_29_48 = multiplicand[19] & multiplier[29];
  assign pp_29_49 = multiplicand[20] & multiplier[29];
  assign pp_29_50 = multiplicand[21] & multiplier[29];
  assign pp_29_51 = multiplicand[22] & multiplier[29];
  assign pp_29_52 = multiplicand[23] & multiplier[29];
  assign pp_29_53 = multiplicand[24] & multiplier[29];
  assign pp_29_54 = multiplicand[25] & multiplier[29];
  assign pp_29_55 = multiplicand[26] & multiplier[29];
  assign pp_29_56 = multiplicand[27] & multiplier[29];
  assign pp_29_57 = multiplicand[28] & multiplier[29];
  assign pp_29_58 = multiplicand[29] & multiplier[29];
  assign pp_29_59 = multiplicand[30] & multiplier[29];
  assign pp_29_60 = multiplicand[31] & multiplier[29];
  assign pp_2_10 = multiplicand[8] & multiplier[2];
  assign pp_2_11 = multiplicand[9] & multiplier[2];
  assign pp_2_12 = multiplicand[10] & multiplier[2];
  assign pp_2_13 = multiplicand[11] & multiplier[2];
  assign pp_2_14 = multiplicand[12] & multiplier[2];
  assign pp_2_15 = multiplicand[13] & multiplier[2];
  assign pp_2_16 = multiplicand[14] & multiplier[2];
  assign pp_2_17 = multiplicand[15] & multiplier[2];
  assign pp_2_18 = multiplicand[16] & multiplier[2];
  assign pp_2_19 = multiplicand[17] & multiplier[2];
  assign pp_2_2 = multiplicand[0] & multiplier[2];
  assign pp_2_20 = multiplicand[18] & multiplier[2];
  assign pp_2_21 = multiplicand[19] & multiplier[2];
  assign pp_2_22 = multiplicand[20] & multiplier[2];
  assign pp_2_23 = multiplicand[21] & multiplier[2];
  assign pp_2_24 = multiplicand[22] & multiplier[2];
  assign pp_2_25 = multiplicand[23] & multiplier[2];
  assign pp_2_26 = multiplicand[24] & multiplier[2];
  assign pp_2_27 = multiplicand[25] & multiplier[2];
  assign pp_2_28 = multiplicand[26] & multiplier[2];
  assign pp_2_29 = multiplicand[27] & multiplier[2];
  assign pp_2_3 = multiplicand[1] & multiplier[2];
  assign pp_2_30 = multiplicand[28] & multiplier[2];
  assign pp_2_31 = multiplicand[29] & multiplier[2];
  assign pp_2_32 = multiplicand[30] & multiplier[2];
  assign pp_2_33 = multiplicand[31] & multiplier[2];
  assign pp_2_4 = multiplicand[2] & multiplier[2];
  assign pp_2_5 = multiplicand[3] & multiplier[2];
  assign pp_2_6 = multiplicand[4] & multiplier[2];
  assign pp_2_7 = multiplicand[5] & multiplier[2];
  assign pp_2_8 = multiplicand[6] & multiplier[2];
  assign pp_2_9 = multiplicand[7] & multiplier[2];
  assign pp_30_30 = multiplicand[0] & multiplier[30];
  assign pp_30_31 = multiplicand[1] & multiplier[30];
  assign pp_30_32 = multiplicand[2] & multiplier[30];
  assign pp_30_33 = multiplicand[3] & multiplier[30];
  assign pp_30_34 = multiplicand[4] & multiplier[30];
  assign pp_30_35 = multiplicand[5] & multiplier[30];
  assign pp_30_36 = multiplicand[6] & multiplier[30];
  assign pp_30_37 = multiplicand[7] & multiplier[30];
  assign pp_30_38 = multiplicand[8] & multiplier[30];
  assign pp_30_39 = multiplicand[9] & multiplier[30];
  assign pp_30_40 = multiplicand[10] & multiplier[30];
  assign pp_30_41 = multiplicand[11] & multiplier[30];
  assign pp_30_42 = multiplicand[12] & multiplier[30];
  assign pp_30_43 = multiplicand[13] & multiplier[30];
  assign pp_30_44 = multiplicand[14] & multiplier[30];
  assign pp_30_45 = multiplicand[15] & multiplier[30];
  assign pp_30_46 = multiplicand[16] & multiplier[30];
  assign pp_30_47 = multiplicand[17] & multiplier[30];
  assign pp_30_48 = multiplicand[18] & multiplier[30];
  assign pp_30_49 = multiplicand[19] & multiplier[30];
  assign pp_30_50 = multiplicand[20] & multiplier[30];
  assign pp_30_51 = multiplicand[21] & multiplier[30];
  assign pp_30_52 = multiplicand[22] & multiplier[30];
  assign pp_30_53 = multiplicand[23] & multiplier[30];
  assign pp_30_54 = multiplicand[24] & multiplier[30];
  assign pp_30_55 = multiplicand[25] & multiplier[30];
  assign pp_30_56 = multiplicand[26] & multiplier[30];
  assign pp_30_57 = multiplicand[27] & multiplier[30];
  assign pp_30_58 = multiplicand[28] & multiplier[30];
  assign pp_30_59 = multiplicand[29] & multiplier[30];
  assign pp_30_60 = multiplicand[30] & multiplier[30];
  assign pp_30_61 = multiplicand[31] & multiplier[30];
  assign pp_31_31 = multiplicand[0] & multiplier[31];
  assign pp_31_32 = multiplicand[1] & multiplier[31];
  assign pp_31_33 = multiplicand[2] & multiplier[31];
  assign pp_31_34 = multiplicand[3] & multiplier[31];
  assign pp_31_35 = multiplicand[4] & multiplier[31];
  assign pp_31_36 = multiplicand[5] & multiplier[31];
  assign pp_31_37 = multiplicand[6] & multiplier[31];
  assign pp_31_38 = multiplicand[7] & multiplier[31];
  assign pp_31_39 = multiplicand[8] & multiplier[31];
  assign pp_31_40 = multiplicand[9] & multiplier[31];
  assign pp_31_41 = multiplicand[10] & multiplier[31];
  assign pp_31_42 = multiplicand[11] & multiplier[31];
  assign pp_31_43 = multiplicand[12] & multiplier[31];
  assign pp_31_44 = multiplicand[13] & multiplier[31];
  assign pp_31_45 = multiplicand[14] & multiplier[31];
  assign pp_31_46 = multiplicand[15] & multiplier[31];
  assign pp_31_47 = multiplicand[16] & multiplier[31];
  assign pp_31_48 = multiplicand[17] & multiplier[31];
  assign pp_31_49 = multiplicand[18] & multiplier[31];
  assign pp_31_50 = multiplicand[19] & multiplier[31];
  assign pp_31_51 = multiplicand[20] & multiplier[31];
  assign pp_31_52 = multiplicand[21] & multiplier[31];
  assign pp_31_53 = multiplicand[22] & multiplier[31];
  assign pp_31_54 = multiplicand[23] & multiplier[31];
  assign pp_31_55 = multiplicand[24] & multiplier[31];
  assign pp_31_56 = multiplicand[25] & multiplier[31];
  assign pp_31_57 = multiplicand[26] & multiplier[31];
  assign pp_31_58 = multiplicand[27] & multiplier[31];
  assign pp_31_59 = multiplicand[28] & multiplier[31];
  assign pp_31_60 = multiplicand[29] & multiplier[31];
  assign pp_31_61 = multiplicand[30] & multiplier[31];
  assign pp_31_62 = multiplicand[31] & multiplier[31];
  assign pp_3_10 = multiplicand[7] & multiplier[3];
  assign pp_3_11 = multiplicand[8] & multiplier[3];
  assign pp_3_12 = multiplicand[9] & multiplier[3];
  assign pp_3_13 = multiplicand[10] & multiplier[3];
  assign pp_3_14 = multiplicand[11] & multiplier[3];
  assign pp_3_15 = multiplicand[12] & multiplier[3];
  assign pp_3_16 = multiplicand[13] & multiplier[3];
  assign pp_3_17 = multiplicand[14] & multiplier[3];
  assign pp_3_18 = multiplicand[15] & multiplier[3];
  assign pp_3_19 = multiplicand[16] & multiplier[3];
  assign pp_3_20 = multiplicand[17] & multiplier[3];
  assign pp_3_21 = multiplicand[18] & multiplier[3];
  assign pp_3_22 = multiplicand[19] & multiplier[3];
  assign pp_3_23 = multiplicand[20] & multiplier[3];
  assign pp_3_24 = multiplicand[21] & multiplier[3];
  assign pp_3_25 = multiplicand[22] & multiplier[3];
  assign pp_3_26 = multiplicand[23] & multiplier[3];
  assign pp_3_27 = multiplicand[24] & multiplier[3];
  assign pp_3_28 = multiplicand[25] & multiplier[3];
  assign pp_3_29 = multiplicand[26] & multiplier[3];
  assign pp_3_3 = multiplicand[0] & multiplier[3];
  assign pp_3_30 = multiplicand[27] & multiplier[3];
  assign pp_3_31 = multiplicand[28] & multiplier[3];
  assign pp_3_32 = multiplicand[29] & multiplier[3];
  assign pp_3_33 = multiplicand[30] & multiplier[3];
  assign pp_3_34 = multiplicand[31] & multiplier[3];
  assign pp_3_4 = multiplicand[1] & multiplier[3];
  assign pp_3_5 = multiplicand[2] & multiplier[3];
  assign pp_3_6 = multiplicand[3] & multiplier[3];
  assign pp_3_7 = multiplicand[4] & multiplier[3];
  assign pp_3_8 = multiplicand[5] & multiplier[3];
  assign pp_3_9 = multiplicand[6] & multiplier[3];
  assign pp_4_10 = multiplicand[6] & multiplier[4];
  assign pp_4_11 = multiplicand[7] & multiplier[4];
  assign pp_4_12 = multiplicand[8] & multiplier[4];
  assign pp_4_13 = multiplicand[9] & multiplier[4];
  assign pp_4_14 = multiplicand[10] & multiplier[4];
  assign pp_4_15 = multiplicand[11] & multiplier[4];
  assign pp_4_16 = multiplicand[12] & multiplier[4];
  assign pp_4_17 = multiplicand[13] & multiplier[4];
  assign pp_4_18 = multiplicand[14] & multiplier[4];
  assign pp_4_19 = multiplicand[15] & multiplier[4];
  assign pp_4_20 = multiplicand[16] & multiplier[4];
  assign pp_4_21 = multiplicand[17] & multiplier[4];
  assign pp_4_22 = multiplicand[18] & multiplier[4];
  assign pp_4_23 = multiplicand[19] & multiplier[4];
  assign pp_4_24 = multiplicand[20] & multiplier[4];
  assign pp_4_25 = multiplicand[21] & multiplier[4];
  assign pp_4_26 = multiplicand[22] & multiplier[4];
  assign pp_4_27 = multiplicand[23] & multiplier[4];
  assign pp_4_28 = multiplicand[24] & multiplier[4];
  assign pp_4_29 = multiplicand[25] & multiplier[4];
  assign pp_4_30 = multiplicand[26] & multiplier[4];
  assign pp_4_31 = multiplicand[27] & multiplier[4];
  assign pp_4_32 = multiplicand[28] & multiplier[4];
  assign pp_4_33 = multiplicand[29] & multiplier[4];
  assign pp_4_34 = multiplicand[30] & multiplier[4];
  assign pp_4_35 = multiplicand[31] & multiplier[4];
  assign pp_4_4 = multiplicand[0] & multiplier[4];
  assign pp_4_5 = multiplicand[1] & multiplier[4];
  assign pp_4_6 = multiplicand[2] & multiplier[4];
  assign pp_4_7 = multiplicand[3] & multiplier[4];
  assign pp_4_8 = multiplicand[4] & multiplier[4];
  assign pp_4_9 = multiplicand[5] & multiplier[4];
  assign pp_5_10 = multiplicand[5] & multiplier[5];
  assign pp_5_11 = multiplicand[6] & multiplier[5];
  assign pp_5_12 = multiplicand[7] & multiplier[5];
  assign pp_5_13 = multiplicand[8] & multiplier[5];
  assign pp_5_14 = multiplicand[9] & multiplier[5];
  assign pp_5_15 = multiplicand[10] & multiplier[5];
  assign pp_5_16 = multiplicand[11] & multiplier[5];
  assign pp_5_17 = multiplicand[12] & multiplier[5];
  assign pp_5_18 = multiplicand[13] & multiplier[5];
  assign pp_5_19 = multiplicand[14] & multiplier[5];
  assign pp_5_20 = multiplicand[15] & multiplier[5];
  assign pp_5_21 = multiplicand[16] & multiplier[5];
  assign pp_5_22 = multiplicand[17] & multiplier[5];
  assign pp_5_23 = multiplicand[18] & multiplier[5];
  assign pp_5_24 = multiplicand[19] & multiplier[5];
  assign pp_5_25 = multiplicand[20] & multiplier[5];
  assign pp_5_26 = multiplicand[21] & multiplier[5];
  assign pp_5_27 = multiplicand[22] & multiplier[5];
  assign pp_5_28 = multiplicand[23] & multiplier[5];
  assign pp_5_29 = multiplicand[24] & multiplier[5];
  assign pp_5_30 = multiplicand[25] & multiplier[5];
  assign pp_5_31 = multiplicand[26] & multiplier[5];
  assign pp_5_32 = multiplicand[27] & multiplier[5];
  assign pp_5_33 = multiplicand[28] & multiplier[5];
  assign pp_5_34 = multiplicand[29] & multiplier[5];
  assign pp_5_35 = multiplicand[30] & multiplier[5];
  assign pp_5_36 = multiplicand[31] & multiplier[5];
  assign pp_5_5 = multiplicand[0] & multiplier[5];
  assign pp_5_6 = multiplicand[1] & multiplier[5];
  assign pp_5_7 = multiplicand[2] & multiplier[5];
  assign pp_5_8 = multiplicand[3] & multiplier[5];
  assign pp_5_9 = multiplicand[4] & multiplier[5];
  assign pp_6_10 = multiplicand[4] & multiplier[6];
  assign pp_6_11 = multiplicand[5] & multiplier[6];
  assign pp_6_12 = multiplicand[6] & multiplier[6];
  assign pp_6_13 = multiplicand[7] & multiplier[6];
  assign pp_6_14 = multiplicand[8] & multiplier[6];
  assign pp_6_15 = multiplicand[9] & multiplier[6];
  assign pp_6_16 = multiplicand[10] & multiplier[6];
  assign pp_6_17 = multiplicand[11] & multiplier[6];
  assign pp_6_18 = multiplicand[12] & multiplier[6];
  assign pp_6_19 = multiplicand[13] & multiplier[6];
  assign pp_6_20 = multiplicand[14] & multiplier[6];
  assign pp_6_21 = multiplicand[15] & multiplier[6];
  assign pp_6_22 = multiplicand[16] & multiplier[6];
  assign pp_6_23 = multiplicand[17] & multiplier[6];
  assign pp_6_24 = multiplicand[18] & multiplier[6];
  assign pp_6_25 = multiplicand[19] & multiplier[6];
  assign pp_6_26 = multiplicand[20] & multiplier[6];
  assign pp_6_27 = multiplicand[21] & multiplier[6];
  assign pp_6_28 = multiplicand[22] & multiplier[6];
  assign pp_6_29 = multiplicand[23] & multiplier[6];
  assign pp_6_30 = multiplicand[24] & multiplier[6];
  assign pp_6_31 = multiplicand[25] & multiplier[6];
  assign pp_6_32 = multiplicand[26] & multiplier[6];
  assign pp_6_33 = multiplicand[27] & multiplier[6];
  assign pp_6_34 = multiplicand[28] & multiplier[6];
  assign pp_6_35 = multiplicand[29] & multiplier[6];
  assign pp_6_36 = multiplicand[30] & multiplier[6];
  assign pp_6_37 = multiplicand[31] & multiplier[6];
  assign pp_6_6 = multiplicand[0] & multiplier[6];
  assign pp_6_7 = multiplicand[1] & multiplier[6];
  assign pp_6_8 = multiplicand[2] & multiplier[6];
  assign pp_6_9 = multiplicand[3] & multiplier[6];
  assign pp_7_10 = multiplicand[3] & multiplier[7];
  assign pp_7_11 = multiplicand[4] & multiplier[7];
  assign pp_7_12 = multiplicand[5] & multiplier[7];
  assign pp_7_13 = multiplicand[6] & multiplier[7];
  assign pp_7_14 = multiplicand[7] & multiplier[7];
  assign pp_7_15 = multiplicand[8] & multiplier[7];
  assign pp_7_16 = multiplicand[9] & multiplier[7];
  assign pp_7_17 = multiplicand[10] & multiplier[7];
  assign pp_7_18 = multiplicand[11] & multiplier[7];
  assign pp_7_19 = multiplicand[12] & multiplier[7];
  assign pp_7_20 = multiplicand[13] & multiplier[7];
  assign pp_7_21 = multiplicand[14] & multiplier[7];
  assign pp_7_22 = multiplicand[15] & multiplier[7];
  assign pp_7_23 = multiplicand[16] & multiplier[7];
  assign pp_7_24 = multiplicand[17] & multiplier[7];
  assign pp_7_25 = multiplicand[18] & multiplier[7];
  assign pp_7_26 = multiplicand[19] & multiplier[7];
  assign pp_7_27 = multiplicand[20] & multiplier[7];
  assign pp_7_28 = multiplicand[21] & multiplier[7];
  assign pp_7_29 = multiplicand[22] & multiplier[7];
  assign pp_7_30 = multiplicand[23] & multiplier[7];
  assign pp_7_31 = multiplicand[24] & multiplier[7];
  assign pp_7_32 = multiplicand[25] & multiplier[7];
  assign pp_7_33 = multiplicand[26] & multiplier[7];
  assign pp_7_34 = multiplicand[27] & multiplier[7];
  assign pp_7_35 = multiplicand[28] & multiplier[7];
  assign pp_7_36 = multiplicand[29] & multiplier[7];
  assign pp_7_37 = multiplicand[30] & multiplier[7];
  assign pp_7_38 = multiplicand[31] & multiplier[7];
  assign pp_7_7 = multiplicand[0] & multiplier[7];
  assign pp_7_8 = multiplicand[1] & multiplier[7];
  assign pp_7_9 = multiplicand[2] & multiplier[7];
  assign pp_8_10 = multiplicand[2] & multiplier[8];
  assign pp_8_11 = multiplicand[3] & multiplier[8];
  assign pp_8_12 = multiplicand[4] & multiplier[8];
  assign pp_8_13 = multiplicand[5] & multiplier[8];
  assign pp_8_14 = multiplicand[6] & multiplier[8];
  assign pp_8_15 = multiplicand[7] & multiplier[8];
  assign pp_8_16 = multiplicand[8] & multiplier[8];
  assign pp_8_17 = multiplicand[9] & multiplier[8];
  assign pp_8_18 = multiplicand[10] & multiplier[8];
  assign pp_8_19 = multiplicand[11] & multiplier[8];
  assign pp_8_20 = multiplicand[12] & multiplier[8];
  assign pp_8_21 = multiplicand[13] & multiplier[8];
  assign pp_8_22 = multiplicand[14] & multiplier[8];
  assign pp_8_23 = multiplicand[15] & multiplier[8];
  assign pp_8_24 = multiplicand[16] & multiplier[8];
  assign pp_8_25 = multiplicand[17] & multiplier[8];
  assign pp_8_26 = multiplicand[18] & multiplier[8];
  assign pp_8_27 = multiplicand[19] & multiplier[8];
  assign pp_8_28 = multiplicand[20] & multiplier[8];
  assign pp_8_29 = multiplicand[21] & multiplier[8];
  assign pp_8_30 = multiplicand[22] & multiplier[8];
  assign pp_8_31 = multiplicand[23] & multiplier[8];
  assign pp_8_32 = multiplicand[24] & multiplier[8];
  assign pp_8_33 = multiplicand[25] & multiplier[8];
  assign pp_8_34 = multiplicand[26] & multiplier[8];
  assign pp_8_35 = multiplicand[27] & multiplier[8];
  assign pp_8_36 = multiplicand[28] & multiplier[8];
  assign pp_8_37 = multiplicand[29] & multiplier[8];
  assign pp_8_38 = multiplicand[30] & multiplier[8];
  assign pp_8_39 = multiplicand[31] & multiplier[8];
  assign pp_8_8 = multiplicand[0] & multiplier[8];
  assign pp_8_9 = multiplicand[1] & multiplier[8];
  assign pp_9_10 = multiplicand[1] & multiplier[9];
  assign pp_9_11 = multiplicand[2] & multiplier[9];
  assign pp_9_12 = multiplicand[3] & multiplier[9];
  assign pp_9_13 = multiplicand[4] & multiplier[9];
  assign pp_9_14 = multiplicand[5] & multiplier[9];
  assign pp_9_15 = multiplicand[6] & multiplier[9];
  assign pp_9_16 = multiplicand[7] & multiplier[9];
  assign pp_9_17 = multiplicand[8] & multiplier[9];
  assign pp_9_18 = multiplicand[9] & multiplier[9];
  assign pp_9_19 = multiplicand[10] & multiplier[9];
  assign pp_9_20 = multiplicand[11] & multiplier[9];
  assign pp_9_21 = multiplicand[12] & multiplier[9];
  assign pp_9_22 = multiplicand[13] & multiplier[9];
  assign pp_9_23 = multiplicand[14] & multiplier[9];
  assign pp_9_24 = multiplicand[15] & multiplier[9];
  assign pp_9_25 = multiplicand[16] & multiplier[9];
  assign pp_9_26 = multiplicand[17] & multiplier[9];
  assign pp_9_27 = multiplicand[18] & multiplier[9];
  assign pp_9_28 = multiplicand[19] & multiplier[9];
  assign pp_9_29 = multiplicand[20] & multiplier[9];
  assign pp_9_30 = multiplicand[21] & multiplier[9];
  assign pp_9_31 = multiplicand[22] & multiplier[9];
  assign pp_9_32 = multiplicand[23] & multiplier[9];
  assign pp_9_33 = multiplicand[24] & multiplier[9];
  assign pp_9_34 = multiplicand[25] & multiplier[9];
  assign pp_9_35 = multiplicand[26] & multiplier[9];
  assign pp_9_36 = multiplicand[27] & multiplier[9];
  assign pp_9_37 = multiplicand[28] & multiplier[9];
  assign pp_9_38 = multiplicand[29] & multiplier[9];
  assign pp_9_39 = multiplicand[30] & multiplier[9];
  assign pp_9_40 = multiplicand[31] & multiplier[9];
  assign pp_9_9 = multiplicand[0] & multiplier[9];
  wire pp_0_0_0;
  wire pp_0_1_0;
  wire pp_0_1_1;
  wire pp_0_2_0;
  wire pp_0_2_1;
  wire pp_0_2_2;
  wire pp_0_3_0;
  wire pp_0_3_1;
  wire pp_0_3_2;
  wire pp_0_3_3;
  wire pp_0_4_0;
  wire pp_0_4_1;
  wire pp_0_4_2;
  wire pp_0_4_3;
  wire pp_0_4_4;
  wire pp_0_5_0;
  wire pp_0_5_1;
  wire pp_0_5_2;
  wire pp_0_5_3;
  wire pp_0_5_4;
  wire pp_0_5_5;
  wire pp_0_6_0;
  wire pp_0_6_1;
  wire pp_0_6_2;
  wire pp_0_6_3;
  wire pp_0_6_4;
  wire pp_0_6_5;
  wire pp_0_6_6;
  wire pp_0_7_0;
  wire pp_0_7_1;
  wire pp_0_7_2;
  wire pp_0_7_3;
  wire pp_0_7_4;
  wire pp_0_7_5;
  wire pp_0_7_6;
  wire pp_0_7_7;
  wire pp_0_8_0;
  wire pp_0_8_1;
  wire pp_0_8_2;
  wire pp_0_8_3;
  wire pp_0_8_4;
  wire pp_0_8_5;
  wire pp_0_8_6;
  wire pp_0_8_7;
  wire pp_0_8_8;
  wire pp_0_9_0;
  wire pp_0_9_1;
  wire pp_0_9_2;
  wire pp_0_9_3;
  wire pp_0_9_4;
  wire pp_0_9_5;
  wire pp_0_9_6;
  wire pp_0_9_7;
  wire pp_0_9_8;
  wire pp_0_9_9;
  wire pp_0_10_0;
  wire pp_0_10_1;
  wire pp_0_10_2;
  wire pp_0_10_3;
  wire pp_0_10_4;
  wire pp_0_10_5;
  wire pp_0_10_6;
  wire pp_0_10_7;
  wire pp_0_10_8;
  wire pp_0_10_9;
  wire pp_0_10_10;
  wire pp_0_11_0;
  wire pp_0_11_1;
  wire pp_0_11_2;
  wire pp_0_11_3;
  wire pp_0_11_4;
  wire pp_0_11_5;
  wire pp_0_11_6;
  wire pp_0_11_7;
  wire pp_0_11_8;
  wire pp_0_11_9;
  wire pp_0_11_10;
  wire pp_0_11_11;
  wire pp_0_12_0;
  wire pp_0_12_1;
  wire pp_0_12_2;
  wire pp_0_12_3;
  wire pp_0_12_4;
  wire pp_0_12_5;
  wire pp_0_12_6;
  wire pp_0_12_7;
  wire pp_0_12_8;
  wire pp_0_12_9;
  wire pp_0_12_10;
  wire pp_0_12_11;
  wire pp_0_12_12;
  wire pp_0_13_0;
  wire pp_0_13_1;
  wire pp_0_13_2;
  wire pp_0_13_3;
  wire pp_0_13_4;
  wire pp_0_13_5;
  wire pp_0_13_6;
  wire pp_0_13_7;
  wire pp_0_13_8;
  wire pp_0_13_9;
  wire pp_0_13_10;
  wire pp_0_13_11;
  wire pp_0_13_12;
  wire pp_0_13_13;
  wire pp_0_14_0;
  wire pp_0_14_1;
  wire pp_0_14_2;
  wire pp_0_14_3;
  wire pp_0_14_4;
  wire pp_0_14_5;
  wire pp_0_14_6;
  wire pp_0_14_7;
  wire pp_0_14_8;
  wire pp_0_14_9;
  wire pp_0_14_10;
  wire pp_0_14_11;
  wire pp_0_14_12;
  wire pp_0_14_13;
  wire pp_0_14_14;
  wire pp_0_15_0;
  wire pp_0_15_1;
  wire pp_0_15_2;
  wire pp_0_15_3;
  wire pp_0_15_4;
  wire pp_0_15_5;
  wire pp_0_15_6;
  wire pp_0_15_7;
  wire pp_0_15_8;
  wire pp_0_15_9;
  wire pp_0_15_10;
  wire pp_0_15_11;
  wire pp_0_15_12;
  wire pp_0_15_13;
  wire pp_0_15_14;
  wire pp_0_15_15;
  wire pp_0_16_0;
  wire pp_0_16_1;
  wire pp_0_16_2;
  wire pp_0_16_3;
  wire pp_0_16_4;
  wire pp_0_16_5;
  wire pp_0_16_6;
  wire pp_0_16_7;
  wire pp_0_16_8;
  wire pp_0_16_9;
  wire pp_0_16_10;
  wire pp_0_16_11;
  wire pp_0_16_12;
  wire pp_0_16_13;
  wire pp_0_16_14;
  wire pp_0_16_15;
  wire pp_0_16_16;
  wire pp_0_17_0;
  wire pp_0_17_1;
  wire pp_0_17_2;
  wire pp_0_17_3;
  wire pp_0_17_4;
  wire pp_0_17_5;
  wire pp_0_17_6;
  wire pp_0_17_7;
  wire pp_0_17_8;
  wire pp_0_17_9;
  wire pp_0_17_10;
  wire pp_0_17_11;
  wire pp_0_17_12;
  wire pp_0_17_13;
  wire pp_0_17_14;
  wire pp_0_17_15;
  wire pp_0_17_16;
  wire pp_0_17_17;
  wire pp_0_18_0;
  wire pp_0_18_1;
  wire pp_0_18_2;
  wire pp_0_18_3;
  wire pp_0_18_4;
  wire pp_0_18_5;
  wire pp_0_18_6;
  wire pp_0_18_7;
  wire pp_0_18_8;
  wire pp_0_18_9;
  wire pp_0_18_10;
  wire pp_0_18_11;
  wire pp_0_18_12;
  wire pp_0_18_13;
  wire pp_0_18_14;
  wire pp_0_18_15;
  wire pp_0_18_16;
  wire pp_0_18_17;
  wire pp_0_18_18;
  wire pp_0_19_0;
  wire pp_0_19_1;
  wire pp_0_19_2;
  wire pp_0_19_3;
  wire pp_0_19_4;
  wire pp_0_19_5;
  wire pp_0_19_6;
  wire pp_0_19_7;
  wire pp_0_19_8;
  wire pp_0_19_9;
  wire pp_0_19_10;
  wire pp_0_19_11;
  wire pp_0_19_12;
  wire pp_0_19_13;
  wire pp_0_19_14;
  wire pp_0_19_15;
  wire pp_0_19_16;
  wire pp_0_19_17;
  wire pp_0_19_18;
  wire pp_0_19_19;
  wire pp_0_20_0;
  wire pp_0_20_1;
  wire pp_0_20_2;
  wire pp_0_20_3;
  wire pp_0_20_4;
  wire pp_0_20_5;
  wire pp_0_20_6;
  wire pp_0_20_7;
  wire pp_0_20_8;
  wire pp_0_20_9;
  wire pp_0_20_10;
  wire pp_0_20_11;
  wire pp_0_20_12;
  wire pp_0_20_13;
  wire pp_0_20_14;
  wire pp_0_20_15;
  wire pp_0_20_16;
  wire pp_0_20_17;
  wire pp_0_20_18;
  wire pp_0_20_19;
  wire pp_0_20_20;
  wire pp_0_21_0;
  wire pp_0_21_1;
  wire pp_0_21_2;
  wire pp_0_21_3;
  wire pp_0_21_4;
  wire pp_0_21_5;
  wire pp_0_21_6;
  wire pp_0_21_7;
  wire pp_0_21_8;
  wire pp_0_21_9;
  wire pp_0_21_10;
  wire pp_0_21_11;
  wire pp_0_21_12;
  wire pp_0_21_13;
  wire pp_0_21_14;
  wire pp_0_21_15;
  wire pp_0_21_16;
  wire pp_0_21_17;
  wire pp_0_21_18;
  wire pp_0_21_19;
  wire pp_0_21_20;
  wire pp_0_21_21;
  wire pp_0_22_0;
  wire pp_0_22_1;
  wire pp_0_22_2;
  wire pp_0_22_3;
  wire pp_0_22_4;
  wire pp_0_22_5;
  wire pp_0_22_6;
  wire pp_0_22_7;
  wire pp_0_22_8;
  wire pp_0_22_9;
  wire pp_0_22_10;
  wire pp_0_22_11;
  wire pp_0_22_12;
  wire pp_0_22_13;
  wire pp_0_22_14;
  wire pp_0_22_15;
  wire pp_0_22_16;
  wire pp_0_22_17;
  wire pp_0_22_18;
  wire pp_0_22_19;
  wire pp_0_22_20;
  wire pp_0_22_21;
  wire pp_0_22_22;
  wire pp_0_23_0;
  wire pp_0_23_1;
  wire pp_0_23_2;
  wire pp_0_23_3;
  wire pp_0_23_4;
  wire pp_0_23_5;
  wire pp_0_23_6;
  wire pp_0_23_7;
  wire pp_0_23_8;
  wire pp_0_23_9;
  wire pp_0_23_10;
  wire pp_0_23_11;
  wire pp_0_23_12;
  wire pp_0_23_13;
  wire pp_0_23_14;
  wire pp_0_23_15;
  wire pp_0_23_16;
  wire pp_0_23_17;
  wire pp_0_23_18;
  wire pp_0_23_19;
  wire pp_0_23_20;
  wire pp_0_23_21;
  wire pp_0_23_22;
  wire pp_0_23_23;
  wire pp_0_24_0;
  wire pp_0_24_1;
  wire pp_0_24_2;
  wire pp_0_24_3;
  wire pp_0_24_4;
  wire pp_0_24_5;
  wire pp_0_24_6;
  wire pp_0_24_7;
  wire pp_0_24_8;
  wire pp_0_24_9;
  wire pp_0_24_10;
  wire pp_0_24_11;
  wire pp_0_24_12;
  wire pp_0_24_13;
  wire pp_0_24_14;
  wire pp_0_24_15;
  wire pp_0_24_16;
  wire pp_0_24_17;
  wire pp_0_24_18;
  wire pp_0_24_19;
  wire pp_0_24_20;
  wire pp_0_24_21;
  wire pp_0_24_22;
  wire pp_0_24_23;
  wire pp_0_24_24;
  wire pp_0_25_0;
  wire pp_0_25_1;
  wire pp_0_25_2;
  wire pp_0_25_3;
  wire pp_0_25_4;
  wire pp_0_25_5;
  wire pp_0_25_6;
  wire pp_0_25_7;
  wire pp_0_25_8;
  wire pp_0_25_9;
  wire pp_0_25_10;
  wire pp_0_25_11;
  wire pp_0_25_12;
  wire pp_0_25_13;
  wire pp_0_25_14;
  wire pp_0_25_15;
  wire pp_0_25_16;
  wire pp_0_25_17;
  wire pp_0_25_18;
  wire pp_0_25_19;
  wire pp_0_25_20;
  wire pp_0_25_21;
  wire pp_0_25_22;
  wire pp_0_25_23;
  wire pp_0_25_24;
  wire pp_0_25_25;
  wire pp_0_26_0;
  wire pp_0_26_1;
  wire pp_0_26_2;
  wire pp_0_26_3;
  wire pp_0_26_4;
  wire pp_0_26_5;
  wire pp_0_26_6;
  wire pp_0_26_7;
  wire pp_0_26_8;
  wire pp_0_26_9;
  wire pp_0_26_10;
  wire pp_0_26_11;
  wire pp_0_26_12;
  wire pp_0_26_13;
  wire pp_0_26_14;
  wire pp_0_26_15;
  wire pp_0_26_16;
  wire pp_0_26_17;
  wire pp_0_26_18;
  wire pp_0_26_19;
  wire pp_0_26_20;
  wire pp_0_26_21;
  wire pp_0_26_22;
  wire pp_0_26_23;
  wire pp_0_26_24;
  wire pp_0_26_25;
  wire pp_0_26_26;
  wire pp_0_27_0;
  wire pp_0_27_1;
  wire pp_0_27_2;
  wire pp_0_27_3;
  wire pp_0_27_4;
  wire pp_0_27_5;
  wire pp_0_27_6;
  wire pp_0_27_7;
  wire pp_0_27_8;
  wire pp_0_27_9;
  wire pp_0_27_10;
  wire pp_0_27_11;
  wire pp_0_27_12;
  wire pp_0_27_13;
  wire pp_0_27_14;
  wire pp_0_27_15;
  wire pp_0_27_16;
  wire pp_0_27_17;
  wire pp_0_27_18;
  wire pp_0_27_19;
  wire pp_0_27_20;
  wire pp_0_27_21;
  wire pp_0_27_22;
  wire pp_0_27_23;
  wire pp_0_27_24;
  wire pp_0_27_25;
  wire pp_0_27_26;
  wire pp_0_27_27;
  wire pp_0_28_0;
  wire pp_0_28_1;
  wire pp_0_28_2;
  wire pp_0_28_3;
  wire pp_0_28_4;
  wire pp_0_28_5;
  wire pp_0_28_6;
  wire pp_0_28_7;
  wire pp_0_28_8;
  wire pp_0_28_9;
  wire pp_0_28_10;
  wire pp_0_28_11;
  wire pp_0_28_12;
  wire pp_0_28_13;
  wire pp_0_28_14;
  wire pp_0_28_15;
  wire pp_0_28_16;
  wire pp_0_28_17;
  wire pp_0_28_18;
  wire pp_0_28_19;
  wire pp_0_28_20;
  wire pp_0_28_21;
  wire pp_0_28_22;
  wire pp_0_28_23;
  wire pp_0_28_24;
  wire pp_0_28_25;
  wire pp_0_28_26;
  wire pp_0_28_27;
  wire pp_0_28_28;
  wire pp_0_29_0;
  wire pp_0_29_1;
  wire pp_0_29_2;
  wire pp_0_29_3;
  wire pp_0_29_4;
  wire pp_0_29_5;
  wire pp_0_29_6;
  wire pp_0_29_7;
  wire pp_0_29_8;
  wire pp_0_29_9;
  wire pp_0_29_10;
  wire pp_0_29_11;
  wire pp_0_29_12;
  wire pp_0_29_13;
  wire pp_0_29_14;
  wire pp_0_29_15;
  wire pp_0_29_16;
  wire pp_0_29_17;
  wire pp_0_29_18;
  wire pp_0_29_19;
  wire pp_0_29_20;
  wire pp_0_29_21;
  wire pp_0_29_22;
  wire pp_0_29_23;
  wire pp_0_29_24;
  wire pp_0_29_25;
  wire pp_0_29_26;
  wire pp_0_29_27;
  wire pp_0_29_28;
  wire pp_0_29_29;
  wire pp_0_30_0;
  wire pp_0_30_1;
  wire pp_0_30_2;
  wire pp_0_30_3;
  wire pp_0_30_4;
  wire pp_0_30_5;
  wire pp_0_30_6;
  wire pp_0_30_7;
  wire pp_0_30_8;
  wire pp_0_30_9;
  wire pp_0_30_10;
  wire pp_0_30_11;
  wire pp_0_30_12;
  wire pp_0_30_13;
  wire pp_0_30_14;
  wire pp_0_30_15;
  wire pp_0_30_16;
  wire pp_0_30_17;
  wire pp_0_30_18;
  wire pp_0_30_19;
  wire pp_0_30_20;
  wire pp_0_30_21;
  wire pp_0_30_22;
  wire pp_0_30_23;
  wire pp_0_30_24;
  wire pp_0_30_25;
  wire pp_0_30_26;
  wire pp_0_30_27;
  wire pp_0_30_28;
  wire pp_0_30_29;
  wire pp_0_30_30;
  wire pp_0_31_0;
  wire pp_0_31_1;
  wire pp_0_31_2;
  wire pp_0_31_3;
  wire pp_0_31_4;
  wire pp_0_31_5;
  wire pp_0_31_6;
  wire pp_0_31_7;
  wire pp_0_31_8;
  wire pp_0_31_9;
  wire pp_0_31_10;
  wire pp_0_31_11;
  wire pp_0_31_12;
  wire pp_0_31_13;
  wire pp_0_31_14;
  wire pp_0_31_15;
  wire pp_0_31_16;
  wire pp_0_31_17;
  wire pp_0_31_18;
  wire pp_0_31_19;
  wire pp_0_31_20;
  wire pp_0_31_21;
  wire pp_0_31_22;
  wire pp_0_31_23;
  wire pp_0_31_24;
  wire pp_0_31_25;
  wire pp_0_31_26;
  wire pp_0_31_27;
  wire pp_0_31_28;
  wire pp_0_31_29;
  wire pp_0_31_30;
  wire pp_0_31_31;
  wire pp_0_32_0;
  wire pp_0_32_1;
  wire pp_0_32_2;
  wire pp_0_32_3;
  wire pp_0_32_4;
  wire pp_0_32_5;
  wire pp_0_32_6;
  wire pp_0_32_7;
  wire pp_0_32_8;
  wire pp_0_32_9;
  wire pp_0_32_10;
  wire pp_0_32_11;
  wire pp_0_32_12;
  wire pp_0_32_13;
  wire pp_0_32_14;
  wire pp_0_32_15;
  wire pp_0_32_16;
  wire pp_0_32_17;
  wire pp_0_32_18;
  wire pp_0_32_19;
  wire pp_0_32_20;
  wire pp_0_32_21;
  wire pp_0_32_22;
  wire pp_0_32_23;
  wire pp_0_32_24;
  wire pp_0_32_25;
  wire pp_0_32_26;
  wire pp_0_32_27;
  wire pp_0_32_28;
  wire pp_0_32_29;
  wire pp_0_32_30;
  wire pp_0_33_0;
  wire pp_0_33_1;
  wire pp_0_33_2;
  wire pp_0_33_3;
  wire pp_0_33_4;
  wire pp_0_33_5;
  wire pp_0_33_6;
  wire pp_0_33_7;
  wire pp_0_33_8;
  wire pp_0_33_9;
  wire pp_0_33_10;
  wire pp_0_33_11;
  wire pp_0_33_12;
  wire pp_0_33_13;
  wire pp_0_33_14;
  wire pp_0_33_15;
  wire pp_0_33_16;
  wire pp_0_33_17;
  wire pp_0_33_18;
  wire pp_0_33_19;
  wire pp_0_33_20;
  wire pp_0_33_21;
  wire pp_0_33_22;
  wire pp_0_33_23;
  wire pp_0_33_24;
  wire pp_0_33_25;
  wire pp_0_33_26;
  wire pp_0_33_27;
  wire pp_0_33_28;
  wire pp_0_33_29;
  wire pp_0_34_0;
  wire pp_0_34_1;
  wire pp_0_34_2;
  wire pp_0_34_3;
  wire pp_0_34_4;
  wire pp_0_34_5;
  wire pp_0_34_6;
  wire pp_0_34_7;
  wire pp_0_34_8;
  wire pp_0_34_9;
  wire pp_0_34_10;
  wire pp_0_34_11;
  wire pp_0_34_12;
  wire pp_0_34_13;
  wire pp_0_34_14;
  wire pp_0_34_15;
  wire pp_0_34_16;
  wire pp_0_34_17;
  wire pp_0_34_18;
  wire pp_0_34_19;
  wire pp_0_34_20;
  wire pp_0_34_21;
  wire pp_0_34_22;
  wire pp_0_34_23;
  wire pp_0_34_24;
  wire pp_0_34_25;
  wire pp_0_34_26;
  wire pp_0_34_27;
  wire pp_0_34_28;
  wire pp_0_35_0;
  wire pp_0_35_1;
  wire pp_0_35_2;
  wire pp_0_35_3;
  wire pp_0_35_4;
  wire pp_0_35_5;
  wire pp_0_35_6;
  wire pp_0_35_7;
  wire pp_0_35_8;
  wire pp_0_35_9;
  wire pp_0_35_10;
  wire pp_0_35_11;
  wire pp_0_35_12;
  wire pp_0_35_13;
  wire pp_0_35_14;
  wire pp_0_35_15;
  wire pp_0_35_16;
  wire pp_0_35_17;
  wire pp_0_35_18;
  wire pp_0_35_19;
  wire pp_0_35_20;
  wire pp_0_35_21;
  wire pp_0_35_22;
  wire pp_0_35_23;
  wire pp_0_35_24;
  wire pp_0_35_25;
  wire pp_0_35_26;
  wire pp_0_35_27;
  wire pp_0_36_0;
  wire pp_0_36_1;
  wire pp_0_36_2;
  wire pp_0_36_3;
  wire pp_0_36_4;
  wire pp_0_36_5;
  wire pp_0_36_6;
  wire pp_0_36_7;
  wire pp_0_36_8;
  wire pp_0_36_9;
  wire pp_0_36_10;
  wire pp_0_36_11;
  wire pp_0_36_12;
  wire pp_0_36_13;
  wire pp_0_36_14;
  wire pp_0_36_15;
  wire pp_0_36_16;
  wire pp_0_36_17;
  wire pp_0_36_18;
  wire pp_0_36_19;
  wire pp_0_36_20;
  wire pp_0_36_21;
  wire pp_0_36_22;
  wire pp_0_36_23;
  wire pp_0_36_24;
  wire pp_0_36_25;
  wire pp_0_36_26;
  wire pp_0_37_0;
  wire pp_0_37_1;
  wire pp_0_37_2;
  wire pp_0_37_3;
  wire pp_0_37_4;
  wire pp_0_37_5;
  wire pp_0_37_6;
  wire pp_0_37_7;
  wire pp_0_37_8;
  wire pp_0_37_9;
  wire pp_0_37_10;
  wire pp_0_37_11;
  wire pp_0_37_12;
  wire pp_0_37_13;
  wire pp_0_37_14;
  wire pp_0_37_15;
  wire pp_0_37_16;
  wire pp_0_37_17;
  wire pp_0_37_18;
  wire pp_0_37_19;
  wire pp_0_37_20;
  wire pp_0_37_21;
  wire pp_0_37_22;
  wire pp_0_37_23;
  wire pp_0_37_24;
  wire pp_0_37_25;
  wire pp_0_38_0;
  wire pp_0_38_1;
  wire pp_0_38_2;
  wire pp_0_38_3;
  wire pp_0_38_4;
  wire pp_0_38_5;
  wire pp_0_38_6;
  wire pp_0_38_7;
  wire pp_0_38_8;
  wire pp_0_38_9;
  wire pp_0_38_10;
  wire pp_0_38_11;
  wire pp_0_38_12;
  wire pp_0_38_13;
  wire pp_0_38_14;
  wire pp_0_38_15;
  wire pp_0_38_16;
  wire pp_0_38_17;
  wire pp_0_38_18;
  wire pp_0_38_19;
  wire pp_0_38_20;
  wire pp_0_38_21;
  wire pp_0_38_22;
  wire pp_0_38_23;
  wire pp_0_38_24;
  wire pp_0_39_0;
  wire pp_0_39_1;
  wire pp_0_39_2;
  wire pp_0_39_3;
  wire pp_0_39_4;
  wire pp_0_39_5;
  wire pp_0_39_6;
  wire pp_0_39_7;
  wire pp_0_39_8;
  wire pp_0_39_9;
  wire pp_0_39_10;
  wire pp_0_39_11;
  wire pp_0_39_12;
  wire pp_0_39_13;
  wire pp_0_39_14;
  wire pp_0_39_15;
  wire pp_0_39_16;
  wire pp_0_39_17;
  wire pp_0_39_18;
  wire pp_0_39_19;
  wire pp_0_39_20;
  wire pp_0_39_21;
  wire pp_0_39_22;
  wire pp_0_39_23;
  wire pp_0_40_0;
  wire pp_0_40_1;
  wire pp_0_40_2;
  wire pp_0_40_3;
  wire pp_0_40_4;
  wire pp_0_40_5;
  wire pp_0_40_6;
  wire pp_0_40_7;
  wire pp_0_40_8;
  wire pp_0_40_9;
  wire pp_0_40_10;
  wire pp_0_40_11;
  wire pp_0_40_12;
  wire pp_0_40_13;
  wire pp_0_40_14;
  wire pp_0_40_15;
  wire pp_0_40_16;
  wire pp_0_40_17;
  wire pp_0_40_18;
  wire pp_0_40_19;
  wire pp_0_40_20;
  wire pp_0_40_21;
  wire pp_0_40_22;
  wire pp_0_41_0;
  wire pp_0_41_1;
  wire pp_0_41_2;
  wire pp_0_41_3;
  wire pp_0_41_4;
  wire pp_0_41_5;
  wire pp_0_41_6;
  wire pp_0_41_7;
  wire pp_0_41_8;
  wire pp_0_41_9;
  wire pp_0_41_10;
  wire pp_0_41_11;
  wire pp_0_41_12;
  wire pp_0_41_13;
  wire pp_0_41_14;
  wire pp_0_41_15;
  wire pp_0_41_16;
  wire pp_0_41_17;
  wire pp_0_41_18;
  wire pp_0_41_19;
  wire pp_0_41_20;
  wire pp_0_41_21;
  wire pp_0_42_0;
  wire pp_0_42_1;
  wire pp_0_42_2;
  wire pp_0_42_3;
  wire pp_0_42_4;
  wire pp_0_42_5;
  wire pp_0_42_6;
  wire pp_0_42_7;
  wire pp_0_42_8;
  wire pp_0_42_9;
  wire pp_0_42_10;
  wire pp_0_42_11;
  wire pp_0_42_12;
  wire pp_0_42_13;
  wire pp_0_42_14;
  wire pp_0_42_15;
  wire pp_0_42_16;
  wire pp_0_42_17;
  wire pp_0_42_18;
  wire pp_0_42_19;
  wire pp_0_42_20;
  wire pp_0_43_0;
  wire pp_0_43_1;
  wire pp_0_43_2;
  wire pp_0_43_3;
  wire pp_0_43_4;
  wire pp_0_43_5;
  wire pp_0_43_6;
  wire pp_0_43_7;
  wire pp_0_43_8;
  wire pp_0_43_9;
  wire pp_0_43_10;
  wire pp_0_43_11;
  wire pp_0_43_12;
  wire pp_0_43_13;
  wire pp_0_43_14;
  wire pp_0_43_15;
  wire pp_0_43_16;
  wire pp_0_43_17;
  wire pp_0_43_18;
  wire pp_0_43_19;
  wire pp_0_44_0;
  wire pp_0_44_1;
  wire pp_0_44_2;
  wire pp_0_44_3;
  wire pp_0_44_4;
  wire pp_0_44_5;
  wire pp_0_44_6;
  wire pp_0_44_7;
  wire pp_0_44_8;
  wire pp_0_44_9;
  wire pp_0_44_10;
  wire pp_0_44_11;
  wire pp_0_44_12;
  wire pp_0_44_13;
  wire pp_0_44_14;
  wire pp_0_44_15;
  wire pp_0_44_16;
  wire pp_0_44_17;
  wire pp_0_44_18;
  wire pp_0_45_0;
  wire pp_0_45_1;
  wire pp_0_45_2;
  wire pp_0_45_3;
  wire pp_0_45_4;
  wire pp_0_45_5;
  wire pp_0_45_6;
  wire pp_0_45_7;
  wire pp_0_45_8;
  wire pp_0_45_9;
  wire pp_0_45_10;
  wire pp_0_45_11;
  wire pp_0_45_12;
  wire pp_0_45_13;
  wire pp_0_45_14;
  wire pp_0_45_15;
  wire pp_0_45_16;
  wire pp_0_45_17;
  wire pp_0_46_0;
  wire pp_0_46_1;
  wire pp_0_46_2;
  wire pp_0_46_3;
  wire pp_0_46_4;
  wire pp_0_46_5;
  wire pp_0_46_6;
  wire pp_0_46_7;
  wire pp_0_46_8;
  wire pp_0_46_9;
  wire pp_0_46_10;
  wire pp_0_46_11;
  wire pp_0_46_12;
  wire pp_0_46_13;
  wire pp_0_46_14;
  wire pp_0_46_15;
  wire pp_0_46_16;
  wire pp_0_47_0;
  wire pp_0_47_1;
  wire pp_0_47_2;
  wire pp_0_47_3;
  wire pp_0_47_4;
  wire pp_0_47_5;
  wire pp_0_47_6;
  wire pp_0_47_7;
  wire pp_0_47_8;
  wire pp_0_47_9;
  wire pp_0_47_10;
  wire pp_0_47_11;
  wire pp_0_47_12;
  wire pp_0_47_13;
  wire pp_0_47_14;
  wire pp_0_47_15;
  wire pp_0_48_0;
  wire pp_0_48_1;
  wire pp_0_48_2;
  wire pp_0_48_3;
  wire pp_0_48_4;
  wire pp_0_48_5;
  wire pp_0_48_6;
  wire pp_0_48_7;
  wire pp_0_48_8;
  wire pp_0_48_9;
  wire pp_0_48_10;
  wire pp_0_48_11;
  wire pp_0_48_12;
  wire pp_0_48_13;
  wire pp_0_48_14;
  wire pp_0_49_0;
  wire pp_0_49_1;
  wire pp_0_49_2;
  wire pp_0_49_3;
  wire pp_0_49_4;
  wire pp_0_49_5;
  wire pp_0_49_6;
  wire pp_0_49_7;
  wire pp_0_49_8;
  wire pp_0_49_9;
  wire pp_0_49_10;
  wire pp_0_49_11;
  wire pp_0_49_12;
  wire pp_0_49_13;
  wire pp_0_50_0;
  wire pp_0_50_1;
  wire pp_0_50_2;
  wire pp_0_50_3;
  wire pp_0_50_4;
  wire pp_0_50_5;
  wire pp_0_50_6;
  wire pp_0_50_7;
  wire pp_0_50_8;
  wire pp_0_50_9;
  wire pp_0_50_10;
  wire pp_0_50_11;
  wire pp_0_50_12;
  wire pp_0_51_0;
  wire pp_0_51_1;
  wire pp_0_51_2;
  wire pp_0_51_3;
  wire pp_0_51_4;
  wire pp_0_51_5;
  wire pp_0_51_6;
  wire pp_0_51_7;
  wire pp_0_51_8;
  wire pp_0_51_9;
  wire pp_0_51_10;
  wire pp_0_51_11;
  wire pp_0_52_0;
  wire pp_0_52_1;
  wire pp_0_52_2;
  wire pp_0_52_3;
  wire pp_0_52_4;
  wire pp_0_52_5;
  wire pp_0_52_6;
  wire pp_0_52_7;
  wire pp_0_52_8;
  wire pp_0_52_9;
  wire pp_0_52_10;
  wire pp_0_53_0;
  wire pp_0_53_1;
  wire pp_0_53_2;
  wire pp_0_53_3;
  wire pp_0_53_4;
  wire pp_0_53_5;
  wire pp_0_53_6;
  wire pp_0_53_7;
  wire pp_0_53_8;
  wire pp_0_53_9;
  wire pp_0_54_0;
  wire pp_0_54_1;
  wire pp_0_54_2;
  wire pp_0_54_3;
  wire pp_0_54_4;
  wire pp_0_54_5;
  wire pp_0_54_6;
  wire pp_0_54_7;
  wire pp_0_54_8;
  wire pp_0_55_0;
  wire pp_0_55_1;
  wire pp_0_55_2;
  wire pp_0_55_3;
  wire pp_0_55_4;
  wire pp_0_55_5;
  wire pp_0_55_6;
  wire pp_0_55_7;
  wire pp_0_56_0;
  wire pp_0_56_1;
  wire pp_0_56_2;
  wire pp_0_56_3;
  wire pp_0_56_4;
  wire pp_0_56_5;
  wire pp_0_56_6;
  wire pp_0_57_0;
  wire pp_0_57_1;
  wire pp_0_57_2;
  wire pp_0_57_3;
  wire pp_0_57_4;
  wire pp_0_57_5;
  wire pp_0_58_0;
  wire pp_0_58_1;
  wire pp_0_58_2;
  wire pp_0_58_3;
  wire pp_0_58_4;
  wire pp_0_59_0;
  wire pp_0_59_1;
  wire pp_0_59_2;
  wire pp_0_59_3;
  wire pp_0_60_0;
  wire pp_0_60_1;
  wire pp_0_60_2;
  wire pp_0_61_0;
  wire pp_0_61_1;
  wire pp_0_62_0;
  wire pp_1_0_0;
  wire pp_1_1_0;
  wire pp_1_1_1;
  wire pp_1_2_0;
  wire pp_1_2_1;
  wire pp_1_2_2;
  wire pp_1_3_0;
  wire pp_1_3_1;
  wire pp_1_3_2;
  wire pp_1_3_3;
  wire pp_1_4_0;
  wire pp_1_4_1;
  wire pp_1_4_2;
  wire pp_1_5_0;
  wire pp_1_5_1;
  wire pp_1_5_2;
  wire pp_1_5_3;
  wire pp_1_5_4;
  wire pp_1_5_5;
  wire pp_1_5_6;
  wire pp_1_6_0;
  wire pp_1_6_1;
  wire pp_1_6_2;
  wire pp_1_6_3;
  wire pp_1_6_4;
  wire pp_1_7_0;
  wire pp_1_7_1;
  wire pp_1_7_2;
  wire pp_1_7_3;
  wire pp_1_7_4;
  wire pp_1_8_0;
  wire pp_1_8_1;
  wire pp_1_8_2;
  wire pp_1_8_3;
  wire pp_1_8_4;
  wire pp_1_8_5;
  wire pp_1_8_6;
  wire pp_1_8_7;
  wire pp_1_8_8;
  wire pp_1_8_9;
  wire pp_1_8_10;
  wire pp_1_9_0;
  wire pp_1_9_1;
  wire pp_1_9_2;
  wire pp_1_9_3;
  wire pp_1_9_4;
  wire pp_1_10_0;
  wire pp_1_10_1;
  wire pp_1_10_2;
  wire pp_1_10_3;
  wire pp_1_10_4;
  wire pp_1_10_5;
  wire pp_1_10_6;
  wire pp_1_10_7;
  wire pp_1_11_0;
  wire pp_1_11_1;
  wire pp_1_11_2;
  wire pp_1_11_3;
  wire pp_1_11_4;
  wire pp_1_11_5;
  wire pp_1_11_6;
  wire pp_1_12_0;
  wire pp_1_12_1;
  wire pp_1_12_2;
  wire pp_1_12_3;
  wire pp_1_12_4;
  wire pp_1_12_5;
  wire pp_1_12_6;
  wire pp_1_12_7;
  wire pp_1_12_8;
  wire pp_1_13_0;
  wire pp_1_13_1;
  wire pp_1_13_2;
  wire pp_1_13_3;
  wire pp_1_13_4;
  wire pp_1_13_5;
  wire pp_1_13_6;
  wire pp_1_13_7;
  wire pp_1_13_8;
  wire pp_1_14_0;
  wire pp_1_14_1;
  wire pp_1_14_2;
  wire pp_1_14_3;
  wire pp_1_14_4;
  wire pp_1_14_5;
  wire pp_1_14_6;
  wire pp_1_14_7;
  wire pp_1_14_8;
  wire pp_1_14_9;
  wire pp_1_15_0;
  wire pp_1_15_1;
  wire pp_1_15_2;
  wire pp_1_15_3;
  wire pp_1_15_4;
  wire pp_1_15_5;
  wire pp_1_15_6;
  wire pp_1_15_7;
  wire pp_1_15_8;
  wire pp_1_15_9;
  wire pp_1_15_10;
  wire pp_1_15_11;
  wire pp_1_16_0;
  wire pp_1_16_1;
  wire pp_1_16_2;
  wire pp_1_16_3;
  wire pp_1_16_4;
  wire pp_1_16_5;
  wire pp_1_16_6;
  wire pp_1_16_7;
  wire pp_1_16_8;
  wire pp_1_16_9;
  wire pp_1_16_10;
  wire pp_1_16_11;
  wire pp_1_17_0;
  wire pp_1_17_1;
  wire pp_1_17_2;
  wire pp_1_17_3;
  wire pp_1_17_4;
  wire pp_1_17_5;
  wire pp_1_17_6;
  wire pp_1_17_7;
  wire pp_1_17_8;
  wire pp_1_17_9;
  wire pp_1_17_10;
  wire pp_1_17_11;
  wire pp_1_17_12;
  wire pp_1_18_0;
  wire pp_1_18_1;
  wire pp_1_18_2;
  wire pp_1_18_3;
  wire pp_1_18_4;
  wire pp_1_18_5;
  wire pp_1_18_6;
  wire pp_1_18_7;
  wire pp_1_18_8;
  wire pp_1_18_9;
  wire pp_1_18_10;
  wire pp_1_18_11;
  wire pp_1_19_0;
  wire pp_1_19_1;
  wire pp_1_19_2;
  wire pp_1_19_3;
  wire pp_1_19_4;
  wire pp_1_19_5;
  wire pp_1_19_6;
  wire pp_1_19_7;
  wire pp_1_19_8;
  wire pp_1_19_9;
  wire pp_1_19_10;
  wire pp_1_19_11;
  wire pp_1_19_12;
  wire pp_1_20_0;
  wire pp_1_20_1;
  wire pp_1_20_2;
  wire pp_1_20_3;
  wire pp_1_20_4;
  wire pp_1_20_5;
  wire pp_1_20_6;
  wire pp_1_20_7;
  wire pp_1_20_8;
  wire pp_1_20_9;
  wire pp_1_20_10;
  wire pp_1_20_11;
  wire pp_1_20_12;
  wire pp_1_20_13;
  wire pp_1_20_14;
  wire pp_1_21_0;
  wire pp_1_21_1;
  wire pp_1_21_2;
  wire pp_1_21_3;
  wire pp_1_21_4;
  wire pp_1_21_5;
  wire pp_1_21_6;
  wire pp_1_21_7;
  wire pp_1_21_8;
  wire pp_1_21_9;
  wire pp_1_21_10;
  wire pp_1_21_11;
  wire pp_1_21_12;
  wire pp_1_21_13;
  wire pp_1_21_14;
  wire pp_1_22_0;
  wire pp_1_22_1;
  wire pp_1_22_2;
  wire pp_1_22_3;
  wire pp_1_22_4;
  wire pp_1_22_5;
  wire pp_1_22_6;
  wire pp_1_22_7;
  wire pp_1_22_8;
  wire pp_1_22_9;
  wire pp_1_22_10;
  wire pp_1_22_11;
  wire pp_1_22_12;
  wire pp_1_22_13;
  wire pp_1_22_14;
  wire pp_1_22_15;
  wire pp_1_23_0;
  wire pp_1_23_1;
  wire pp_1_23_2;
  wire pp_1_23_3;
  wire pp_1_23_4;
  wire pp_1_23_5;
  wire pp_1_23_6;
  wire pp_1_23_7;
  wire pp_1_23_8;
  wire pp_1_23_9;
  wire pp_1_23_10;
  wire pp_1_23_11;
  wire pp_1_23_12;
  wire pp_1_23_13;
  wire pp_1_23_14;
  wire pp_1_24_0;
  wire pp_1_24_1;
  wire pp_1_24_2;
  wire pp_1_24_3;
  wire pp_1_24_4;
  wire pp_1_24_5;
  wire pp_1_24_6;
  wire pp_1_24_7;
  wire pp_1_24_8;
  wire pp_1_24_9;
  wire pp_1_24_10;
  wire pp_1_24_11;
  wire pp_1_24_12;
  wire pp_1_24_13;
  wire pp_1_24_14;
  wire pp_1_24_15;
  wire pp_1_24_16;
  wire pp_1_25_0;
  wire pp_1_25_1;
  wire pp_1_25_2;
  wire pp_1_25_3;
  wire pp_1_25_4;
  wire pp_1_25_5;
  wire pp_1_25_6;
  wire pp_1_25_7;
  wire pp_1_25_8;
  wire pp_1_25_9;
  wire pp_1_25_10;
  wire pp_1_25_11;
  wire pp_1_25_12;
  wire pp_1_25_13;
  wire pp_1_25_14;
  wire pp_1_25_15;
  wire pp_1_25_16;
  wire pp_1_25_17;
  wire pp_1_25_18;
  wire pp_1_25_19;
  wire pp_1_25_20;
  wire pp_1_25_21;
  wire pp_1_25_22;
  wire pp_1_25_23;
  wire pp_1_25_24;
  wire pp_1_25_25;
  wire pp_1_25_26;
  wire pp_1_25_27;
  wire pp_1_25_28;
  wire pp_1_25_29;
  wire pp_1_25_30;
  wire pp_1_25_31;
  wire pp_1_25_32;
  wire pp_1_25_33;
  wire pp_1_26_0;
  wire pp_1_26_1;
  wire pp_1_26_2;
  wire pp_1_26_3;
  wire pp_1_26_4;
  wire pp_1_26_5;
  wire pp_1_26_6;
  wire pp_1_26_7;
  wire pp_1_26_8;
  wire pp_1_26_9;
  wire pp_1_26_10;
  wire pp_1_26_11;
  wire pp_1_27_0;
  wire pp_1_27_1;
  wire pp_1_27_2;
  wire pp_1_27_3;
  wire pp_1_27_4;
  wire pp_1_27_5;
  wire pp_1_27_6;
  wire pp_1_27_7;
  wire pp_1_27_8;
  wire pp_1_27_9;
  wire pp_1_27_10;
  wire pp_1_27_11;
  wire pp_1_27_12;
  wire pp_1_27_13;
  wire pp_1_27_14;
  wire pp_1_27_15;
  wire pp_1_27_16;
  wire pp_1_27_17;
  wire pp_1_28_0;
  wire pp_1_28_1;
  wire pp_1_28_2;
  wire pp_1_28_3;
  wire pp_1_28_4;
  wire pp_1_28_5;
  wire pp_1_28_6;
  wire pp_1_28_7;
  wire pp_1_28_8;
  wire pp_1_28_9;
  wire pp_1_28_10;
  wire pp_1_28_11;
  wire pp_1_28_12;
  wire pp_1_28_13;
  wire pp_1_28_14;
  wire pp_1_28_15;
  wire pp_1_28_16;
  wire pp_1_28_17;
  wire pp_1_28_18;
  wire pp_1_28_19;
  wire pp_1_29_0;
  wire pp_1_29_1;
  wire pp_1_29_2;
  wire pp_1_29_3;
  wire pp_1_29_4;
  wire pp_1_29_5;
  wire pp_1_29_6;
  wire pp_1_29_7;
  wire pp_1_29_8;
  wire pp_1_29_9;
  wire pp_1_29_10;
  wire pp_1_29_11;
  wire pp_1_29_12;
  wire pp_1_29_13;
  wire pp_1_29_14;
  wire pp_1_29_15;
  wire pp_1_29_16;
  wire pp_1_29_17;
  wire pp_1_29_18;
  wire pp_1_30_0;
  wire pp_1_30_1;
  wire pp_1_30_2;
  wire pp_1_30_3;
  wire pp_1_30_4;
  wire pp_1_30_5;
  wire pp_1_30_6;
  wire pp_1_30_7;
  wire pp_1_30_8;
  wire pp_1_30_9;
  wire pp_1_30_10;
  wire pp_1_30_11;
  wire pp_1_30_12;
  wire pp_1_30_13;
  wire pp_1_30_14;
  wire pp_1_30_15;
  wire pp_1_30_16;
  wire pp_1_30_17;
  wire pp_1_30_18;
  wire pp_1_30_19;
  wire pp_1_30_20;
  wire pp_1_31_0;
  wire pp_1_31_1;
  wire pp_1_31_2;
  wire pp_1_31_3;
  wire pp_1_31_4;
  wire pp_1_31_5;
  wire pp_1_31_6;
  wire pp_1_31_7;
  wire pp_1_31_8;
  wire pp_1_31_9;
  wire pp_1_31_10;
  wire pp_1_31_11;
  wire pp_1_31_12;
  wire pp_1_31_13;
  wire pp_1_31_14;
  wire pp_1_31_15;
  wire pp_1_31_16;
  wire pp_1_31_17;
  wire pp_1_31_18;
  wire pp_1_31_19;
  wire pp_1_31_20;
  wire pp_1_31_21;
  wire pp_1_32_0;
  wire pp_1_32_1;
  wire pp_1_32_2;
  wire pp_1_32_3;
  wire pp_1_32_4;
  wire pp_1_32_5;
  wire pp_1_32_6;
  wire pp_1_32_7;
  wire pp_1_32_8;
  wire pp_1_32_9;
  wire pp_1_32_10;
  wire pp_1_32_11;
  wire pp_1_32_12;
  wire pp_1_32_13;
  wire pp_1_32_14;
  wire pp_1_32_15;
  wire pp_1_32_16;
  wire pp_1_32_17;
  wire pp_1_32_18;
  wire pp_1_32_19;
  wire pp_1_32_20;
  wire pp_1_33_0;
  wire pp_1_33_1;
  wire pp_1_33_2;
  wire pp_1_33_3;
  wire pp_1_33_4;
  wire pp_1_33_5;
  wire pp_1_33_6;
  wire pp_1_33_7;
  wire pp_1_33_8;
  wire pp_1_33_9;
  wire pp_1_33_10;
  wire pp_1_33_11;
  wire pp_1_33_12;
  wire pp_1_33_13;
  wire pp_1_33_14;
  wire pp_1_33_15;
  wire pp_1_33_16;
  wire pp_1_33_17;
  wire pp_1_33_18;
  wire pp_1_33_19;
  wire pp_1_34_0;
  wire pp_1_34_1;
  wire pp_1_34_2;
  wire pp_1_34_3;
  wire pp_1_34_4;
  wire pp_1_34_5;
  wire pp_1_34_6;
  wire pp_1_34_7;
  wire pp_1_34_8;
  wire pp_1_34_9;
  wire pp_1_34_10;
  wire pp_1_34_11;
  wire pp_1_34_12;
  wire pp_1_34_13;
  wire pp_1_34_14;
  wire pp_1_34_15;
  wire pp_1_34_16;
  wire pp_1_34_17;
  wire pp_1_34_18;
  wire pp_1_34_19;
  wire pp_1_34_20;
  wire pp_1_35_0;
  wire pp_1_35_1;
  wire pp_1_35_2;
  wire pp_1_35_3;
  wire pp_1_35_4;
  wire pp_1_35_5;
  wire pp_1_35_6;
  wire pp_1_35_7;
  wire pp_1_35_8;
  wire pp_1_35_9;
  wire pp_1_35_10;
  wire pp_1_35_11;
  wire pp_1_35_12;
  wire pp_1_35_13;
  wire pp_1_35_14;
  wire pp_1_35_15;
  wire pp_1_35_16;
  wire pp_1_35_17;
  wire pp_1_35_18;
  wire pp_1_36_0;
  wire pp_1_36_1;
  wire pp_1_36_2;
  wire pp_1_36_3;
  wire pp_1_36_4;
  wire pp_1_36_5;
  wire pp_1_36_6;
  wire pp_1_36_7;
  wire pp_1_36_8;
  wire pp_1_36_9;
  wire pp_1_36_10;
  wire pp_1_36_11;
  wire pp_1_36_12;
  wire pp_1_36_13;
  wire pp_1_36_14;
  wire pp_1_36_15;
  wire pp_1_36_16;
  wire pp_1_36_17;
  wire pp_1_37_0;
  wire pp_1_37_1;
  wire pp_1_37_2;
  wire pp_1_37_3;
  wire pp_1_37_4;
  wire pp_1_37_5;
  wire pp_1_37_6;
  wire pp_1_37_7;
  wire pp_1_37_8;
  wire pp_1_37_9;
  wire pp_1_37_10;
  wire pp_1_37_11;
  wire pp_1_37_12;
  wire pp_1_37_13;
  wire pp_1_37_14;
  wire pp_1_37_15;
  wire pp_1_37_16;
  wire pp_1_37_17;
  wire pp_1_37_18;
  wire pp_1_38_0;
  wire pp_1_38_1;
  wire pp_1_38_2;
  wire pp_1_38_3;
  wire pp_1_38_4;
  wire pp_1_38_5;
  wire pp_1_38_6;
  wire pp_1_38_7;
  wire pp_1_38_8;
  wire pp_1_38_9;
  wire pp_1_38_10;
  wire pp_1_38_11;
  wire pp_1_38_12;
  wire pp_1_38_13;
  wire pp_1_38_14;
  wire pp_1_38_15;
  wire pp_1_38_16;
  wire pp_1_39_0;
  wire pp_1_39_1;
  wire pp_1_39_2;
  wire pp_1_39_3;
  wire pp_1_39_4;
  wire pp_1_39_5;
  wire pp_1_39_6;
  wire pp_1_39_7;
  wire pp_1_39_8;
  wire pp_1_39_9;
  wire pp_1_39_10;
  wire pp_1_39_11;
  wire pp_1_39_12;
  wire pp_1_39_13;
  wire pp_1_39_14;
  wire pp_1_39_15;
  wire pp_1_40_0;
  wire pp_1_40_1;
  wire pp_1_40_2;
  wire pp_1_40_3;
  wire pp_1_40_4;
  wire pp_1_40_5;
  wire pp_1_40_6;
  wire pp_1_40_7;
  wire pp_1_40_8;
  wire pp_1_40_9;
  wire pp_1_40_10;
  wire pp_1_40_11;
  wire pp_1_40_12;
  wire pp_1_40_13;
  wire pp_1_40_14;
  wire pp_1_40_15;
  wire pp_1_40_16;
  wire pp_1_40_17;
  wire pp_1_40_18;
  wire pp_1_40_19;
  wire pp_1_40_20;
  wire pp_1_41_0;
  wire pp_1_41_1;
  wire pp_1_41_2;
  wire pp_1_41_3;
  wire pp_1_41_4;
  wire pp_1_41_5;
  wire pp_1_41_6;
  wire pp_1_41_7;
  wire pp_1_41_8;
  wire pp_1_41_9;
  wire pp_1_41_10;
  wire pp_1_41_11;
  wire pp_1_41_12;
  wire pp_1_41_13;
  wire pp_1_41_14;
  wire pp_1_42_0;
  wire pp_1_42_1;
  wire pp_1_42_2;
  wire pp_1_42_3;
  wire pp_1_42_4;
  wire pp_1_42_5;
  wire pp_1_42_6;
  wire pp_1_42_7;
  wire pp_1_42_8;
  wire pp_1_42_9;
  wire pp_1_42_10;
  wire pp_1_42_11;
  wire pp_1_42_12;
  wire pp_1_43_0;
  wire pp_1_43_1;
  wire pp_1_43_2;
  wire pp_1_43_3;
  wire pp_1_43_4;
  wire pp_1_43_5;
  wire pp_1_43_6;
  wire pp_1_43_7;
  wire pp_1_43_8;
  wire pp_1_43_9;
  wire pp_1_43_10;
  wire pp_1_43_11;
  wire pp_1_43_12;
  wire pp_1_43_13;
  wire pp_1_43_14;
  wire pp_1_44_0;
  wire pp_1_44_1;
  wire pp_1_44_2;
  wire pp_1_44_3;
  wire pp_1_44_4;
  wire pp_1_44_5;
  wire pp_1_44_6;
  wire pp_1_44_7;
  wire pp_1_44_8;
  wire pp_1_44_9;
  wire pp_1_44_10;
  wire pp_1_44_11;
  wire pp_1_44_12;
  wire pp_1_44_13;
  wire pp_1_44_14;
  wire pp_1_44_15;
  wire pp_1_44_16;
  wire pp_1_44_17;
  wire pp_1_44_18;
  wire pp_1_44_19;
  wire pp_1_44_20;
  wire pp_1_44_21;
  wire pp_1_44_22;
  wire pp_1_44_23;
  wire pp_1_44_24;
  wire pp_1_45_0;
  wire pp_1_45_1;
  wire pp_1_45_2;
  wire pp_1_45_3;
  wire pp_1_45_4;
  wire pp_1_45_5;
  wire pp_1_46_0;
  wire pp_1_46_1;
  wire pp_1_46_2;
  wire pp_1_46_3;
  wire pp_1_46_4;
  wire pp_1_46_5;
  wire pp_1_46_6;
  wire pp_1_46_7;
  wire pp_1_46_8;
  wire pp_1_46_9;
  wire pp_1_46_10;
  wire pp_1_46_11;
  wire pp_1_46_12;
  wire pp_1_46_13;
  wire pp_1_46_14;
  wire pp_1_47_0;
  wire pp_1_47_1;
  wire pp_1_47_2;
  wire pp_1_47_3;
  wire pp_1_47_4;
  wire pp_1_47_5;
  wire pp_1_47_6;
  wire pp_1_47_7;
  wire pp_1_47_8;
  wire pp_1_47_9;
  wire pp_1_47_10;
  wire pp_1_47_11;
  wire pp_1_48_0;
  wire pp_1_48_1;
  wire pp_1_48_2;
  wire pp_1_48_3;
  wire pp_1_48_4;
  wire pp_1_48_5;
  wire pp_1_48_6;
  wire pp_1_48_7;
  wire pp_1_48_8;
  wire pp_1_49_0;
  wire pp_1_49_1;
  wire pp_1_49_2;
  wire pp_1_49_3;
  wire pp_1_49_4;
  wire pp_1_49_5;
  wire pp_1_49_6;
  wire pp_1_49_7;
  wire pp_1_49_8;
  wire pp_1_49_9;
  wire pp_1_49_10;
  wire pp_1_50_0;
  wire pp_1_50_1;
  wire pp_1_50_2;
  wire pp_1_50_3;
  wire pp_1_50_4;
  wire pp_1_50_5;
  wire pp_1_50_6;
  wire pp_1_50_7;
  wire pp_1_50_8;
  wire pp_1_51_0;
  wire pp_1_51_1;
  wire pp_1_51_2;
  wire pp_1_51_3;
  wire pp_1_51_4;
  wire pp_1_51_5;
  wire pp_1_51_6;
  wire pp_1_51_7;
  wire pp_1_52_0;
  wire pp_1_52_1;
  wire pp_1_52_2;
  wire pp_1_52_3;
  wire pp_1_52_4;
  wire pp_1_52_5;
  wire pp_1_52_6;
  wire pp_1_52_7;
  wire pp_1_52_8;
  wire pp_1_53_0;
  wire pp_1_53_1;
  wire pp_1_53_2;
  wire pp_1_53_3;
  wire pp_1_53_4;
  wire pp_1_53_5;
  wire pp_1_53_6;
  wire pp_1_54_0;
  wire pp_1_54_1;
  wire pp_1_54_2;
  wire pp_1_54_3;
  wire pp_1_54_4;
  wire pp_1_54_5;
  wire pp_1_55_0;
  wire pp_1_55_1;
  wire pp_1_55_2;
  wire pp_1_55_3;
  wire pp_1_55_4;
  wire pp_1_55_5;
  wire pp_1_55_6;
  wire pp_1_56_0;
  wire pp_1_56_1;
  wire pp_1_56_2;
  wire pp_1_56_3;
  wire pp_1_56_4;
  wire pp_1_56_5;
  wire pp_1_56_6;
  wire pp_1_56_7;
  wire pp_1_56_8;
  wire pp_1_57_0;
  wire pp_1_57_1;
  wire pp_1_58_0;
  wire pp_1_58_1;
  wire pp_1_58_2;
  wire pp_1_58_3;
  wire pp_1_58_4;
  wire pp_1_58_5;
  wire pp_1_58_6;
  wire pp_1_59_0;
  wire pp_1_59_1;
  wire pp_1_59_2;
  wire pp_1_59_3;
  wire pp_1_60_0;
  wire pp_1_61_0;
  wire pp_1_61_1;
  wire pp_1_61_2;
  wire pp_1_62_0;
  wire pp_2_0_0;
  wire pp_2_1_0;
  wire pp_2_1_1;
  wire pp_2_2_0;
  wire pp_2_2_1;
  wire pp_2_2_2;
  wire pp_2_3_0;
  wire pp_2_3_1;
  wire pp_2_3_2;
  wire pp_2_3_3;
  wire pp_2_4_0;
  wire pp_2_4_1;
  wire pp_2_4_2;
  wire pp_2_5_0;
  wire pp_2_5_1;
  wire pp_2_5_2;
  wire pp_2_6_0;
  wire pp_2_6_1;
  wire pp_2_6_2;
  wire pp_2_6_3;
  wire pp_2_6_4;
  wire pp_2_6_5;
  wire pp_2_6_6;
  wire pp_2_7_0;
  wire pp_2_7_1;
  wire pp_2_8_0;
  wire pp_2_8_1;
  wire pp_2_8_2;
  wire pp_2_8_3;
  wire pp_2_8_4;
  wire pp_2_8_5;
  wire pp_2_9_0;
  wire pp_2_9_1;
  wire pp_2_9_2;
  wire pp_2_9_3;
  wire pp_2_9_4;
  wire pp_2_9_5;
  wire pp_2_9_6;
  wire pp_2_9_7;
  wire pp_2_9_8;
  wire pp_2_10_0;
  wire pp_2_10_1;
  wire pp_2_10_2;
  wire pp_2_10_3;
  wire pp_2_11_0;
  wire pp_2_11_1;
  wire pp_2_11_2;
  wire pp_2_11_3;
  wire pp_2_11_4;
  wire pp_2_11_5;
  wire pp_2_11_6;
  wire pp_2_11_7;
  wire pp_2_11_8;
  wire pp_2_12_0;
  wire pp_2_12_1;
  wire pp_2_12_2;
  wire pp_2_13_0;
  wire pp_2_13_1;
  wire pp_2_13_2;
  wire pp_2_13_3;
  wire pp_2_13_4;
  wire pp_2_13_5;
  wire pp_2_14_0;
  wire pp_2_14_1;
  wire pp_2_14_2;
  wire pp_2_14_3;
  wire pp_2_14_4;
  wire pp_2_14_5;
  wire pp_2_14_6;
  wire pp_2_14_7;
  wire pp_2_14_8;
  wire pp_2_14_9;
  wire pp_2_14_10;
  wire pp_2_14_11;
  wire pp_2_14_12;
  wire pp_2_15_0;
  wire pp_2_15_1;
  wire pp_2_15_2;
  wire pp_2_15_3;
  wire pp_2_16_0;
  wire pp_2_16_1;
  wire pp_2_16_2;
  wire pp_2_16_3;
  wire pp_2_16_4;
  wire pp_2_16_5;
  wire pp_2_16_6;
  wire pp_2_16_7;
  wire pp_2_17_0;
  wire pp_2_17_1;
  wire pp_2_17_2;
  wire pp_2_17_3;
  wire pp_2_17_4;
  wire pp_2_17_5;
  wire pp_2_17_6;
  wire pp_2_17_7;
  wire pp_2_17_8;
  wire pp_2_18_0;
  wire pp_2_18_1;
  wire pp_2_18_2;
  wire pp_2_18_3;
  wire pp_2_18_4;
  wire pp_2_18_5;
  wire pp_2_18_6;
  wire pp_2_18_7;
  wire pp_2_19_0;
  wire pp_2_19_1;
  wire pp_2_19_2;
  wire pp_2_19_3;
  wire pp_2_19_4;
  wire pp_2_19_5;
  wire pp_2_19_6;
  wire pp_2_19_7;
  wire pp_2_19_8;
  wire pp_2_20_0;
  wire pp_2_20_1;
  wire pp_2_20_2;
  wire pp_2_20_3;
  wire pp_2_20_4;
  wire pp_2_20_5;
  wire pp_2_20_6;
  wire pp_2_20_7;
  wire pp_2_20_8;
  wire pp_2_21_0;
  wire pp_2_21_1;
  wire pp_2_21_2;
  wire pp_2_21_3;
  wire pp_2_21_4;
  wire pp_2_21_5;
  wire pp_2_21_6;
  wire pp_2_21_7;
  wire pp_2_21_8;
  wire pp_2_21_9;
  wire pp_2_22_0;
  wire pp_2_22_1;
  wire pp_2_22_2;
  wire pp_2_22_3;
  wire pp_2_22_4;
  wire pp_2_22_5;
  wire pp_2_22_6;
  wire pp_2_22_7;
  wire pp_2_22_8;
  wire pp_2_22_9;
  wire pp_2_22_10;
  wire pp_2_22_11;
  wire pp_2_22_12;
  wire pp_2_22_13;
  wire pp_2_22_14;
  wire pp_2_22_15;
  wire pp_2_22_16;
  wire pp_2_22_17;
  wire pp_2_22_18;
  wire pp_2_22_19;
  wire pp_2_22_20;
  wire pp_2_23_0;
  wire pp_2_23_1;
  wire pp_2_23_2;
  wire pp_2_23_3;
  wire pp_2_23_4;
  wire pp_2_24_0;
  wire pp_2_24_1;
  wire pp_2_24_2;
  wire pp_2_24_3;
  wire pp_2_24_4;
  wire pp_2_24_5;
  wire pp_2_24_6;
  wire pp_2_24_7;
  wire pp_2_24_8;
  wire pp_2_24_9;
  wire pp_2_24_10;
  wire pp_2_24_11;
  wire pp_2_25_0;
  wire pp_2_25_1;
  wire pp_2_25_2;
  wire pp_2_25_3;
  wire pp_2_25_4;
  wire pp_2_25_5;
  wire pp_2_25_6;
  wire pp_2_25_7;
  wire pp_2_25_8;
  wire pp_2_25_9;
  wire pp_2_25_10;
  wire pp_2_25_11;
  wire pp_2_25_12;
  wire pp_2_25_13;
  wire pp_2_25_14;
  wire pp_2_25_15;
  wire pp_2_25_16;
  wire pp_2_26_0;
  wire pp_2_26_1;
  wire pp_2_26_2;
  wire pp_2_26_3;
  wire pp_2_26_4;
  wire pp_2_26_5;
  wire pp_2_26_6;
  wire pp_2_26_7;
  wire pp_2_26_8;
  wire pp_2_26_9;
  wire pp_2_26_10;
  wire pp_2_26_11;
  wire pp_2_26_12;
  wire pp_2_26_13;
  wire pp_2_26_14;
  wire pp_2_27_0;
  wire pp_2_27_1;
  wire pp_2_27_2;
  wire pp_2_27_3;
  wire pp_2_27_4;
  wire pp_2_27_5;
  wire pp_2_27_6;
  wire pp_2_27_7;
  wire pp_2_27_8;
  wire pp_2_27_9;
  wire pp_2_27_10;
  wire pp_2_27_11;
  wire pp_2_28_0;
  wire pp_2_28_1;
  wire pp_2_28_2;
  wire pp_2_28_3;
  wire pp_2_28_4;
  wire pp_2_28_5;
  wire pp_2_28_6;
  wire pp_2_28_7;
  wire pp_2_28_8;
  wire pp_2_28_9;
  wire pp_2_28_10;
  wire pp_2_28_11;
  wire pp_2_28_12;
  wire pp_2_29_0;
  wire pp_2_29_1;
  wire pp_2_29_2;
  wire pp_2_29_3;
  wire pp_2_29_4;
  wire pp_2_29_5;
  wire pp_2_29_6;
  wire pp_2_29_7;
  wire pp_2_29_8;
  wire pp_2_29_9;
  wire pp_2_29_10;
  wire pp_2_29_11;
  wire pp_2_29_12;
  wire pp_2_30_0;
  wire pp_2_30_1;
  wire pp_2_30_2;
  wire pp_2_30_3;
  wire pp_2_30_4;
  wire pp_2_30_5;
  wire pp_2_30_6;
  wire pp_2_30_7;
  wire pp_2_30_8;
  wire pp_2_30_9;
  wire pp_2_30_10;
  wire pp_2_30_11;
  wire pp_2_30_12;
  wire pp_2_31_0;
  wire pp_2_31_1;
  wire pp_2_31_2;
  wire pp_2_31_3;
  wire pp_2_31_4;
  wire pp_2_31_5;
  wire pp_2_31_6;
  wire pp_2_31_7;
  wire pp_2_31_8;
  wire pp_2_31_9;
  wire pp_2_31_10;
  wire pp_2_31_11;
  wire pp_2_31_12;
  wire pp_2_31_13;
  wire pp_2_31_14;
  wire pp_2_32_0;
  wire pp_2_32_1;
  wire pp_2_32_2;
  wire pp_2_32_3;
  wire pp_2_32_4;
  wire pp_2_32_5;
  wire pp_2_32_6;
  wire pp_2_32_7;
  wire pp_2_32_8;
  wire pp_2_32_9;
  wire pp_2_32_10;
  wire pp_2_32_11;
  wire pp_2_32_12;
  wire pp_2_32_13;
  wire pp_2_33_0;
  wire pp_2_33_1;
  wire pp_2_33_2;
  wire pp_2_33_3;
  wire pp_2_33_4;
  wire pp_2_33_5;
  wire pp_2_33_6;
  wire pp_2_33_7;
  wire pp_2_33_8;
  wire pp_2_33_9;
  wire pp_2_33_10;
  wire pp_2_33_11;
  wire pp_2_33_12;
  wire pp_2_33_13;
  wire pp_2_33_14;
  wire pp_2_34_0;
  wire pp_2_34_1;
  wire pp_2_34_2;
  wire pp_2_34_3;
  wire pp_2_34_4;
  wire pp_2_34_5;
  wire pp_2_34_6;
  wire pp_2_34_7;
  wire pp_2_34_8;
  wire pp_2_34_9;
  wire pp_2_34_10;
  wire pp_2_34_11;
  wire pp_2_34_12;
  wire pp_2_35_0;
  wire pp_2_35_1;
  wire pp_2_35_2;
  wire pp_2_35_3;
  wire pp_2_35_4;
  wire pp_2_35_5;
  wire pp_2_35_6;
  wire pp_2_35_7;
  wire pp_2_35_8;
  wire pp_2_35_9;
  wire pp_2_35_10;
  wire pp_2_35_11;
  wire pp_2_35_12;
  wire pp_2_35_13;
  wire pp_2_36_0;
  wire pp_2_36_1;
  wire pp_2_36_2;
  wire pp_2_36_3;
  wire pp_2_36_4;
  wire pp_2_36_5;
  wire pp_2_36_6;
  wire pp_2_36_7;
  wire pp_2_36_8;
  wire pp_2_36_9;
  wire pp_2_36_10;
  wire pp_2_36_11;
  wire pp_2_37_0;
  wire pp_2_37_1;
  wire pp_2_37_2;
  wire pp_2_37_3;
  wire pp_2_37_4;
  wire pp_2_37_5;
  wire pp_2_37_6;
  wire pp_2_37_7;
  wire pp_2_37_8;
  wire pp_2_37_9;
  wire pp_2_37_10;
  wire pp_2_37_11;
  wire pp_2_37_12;
  wire pp_2_38_0;
  wire pp_2_38_1;
  wire pp_2_38_2;
  wire pp_2_38_3;
  wire pp_2_38_4;
  wire pp_2_38_5;
  wire pp_2_38_6;
  wire pp_2_38_7;
  wire pp_2_38_8;
  wire pp_2_38_9;
  wire pp_2_38_10;
  wire pp_2_38_11;
  wire pp_2_38_12;
  wire pp_2_39_0;
  wire pp_2_39_1;
  wire pp_2_39_2;
  wire pp_2_39_3;
  wire pp_2_39_4;
  wire pp_2_39_5;
  wire pp_2_39_6;
  wire pp_2_39_7;
  wire pp_2_39_8;
  wire pp_2_39_9;
  wire pp_2_39_10;
  wire pp_2_40_0;
  wire pp_2_40_1;
  wire pp_2_40_2;
  wire pp_2_40_3;
  wire pp_2_40_4;
  wire pp_2_40_5;
  wire pp_2_40_6;
  wire pp_2_40_7;
  wire pp_2_40_8;
  wire pp_2_40_9;
  wire pp_2_40_10;
  wire pp_2_40_11;
  wire pp_2_41_0;
  wire pp_2_41_1;
  wire pp_2_41_2;
  wire pp_2_41_3;
  wire pp_2_41_4;
  wire pp_2_41_5;
  wire pp_2_41_6;
  wire pp_2_41_7;
  wire pp_2_41_8;
  wire pp_2_41_9;
  wire pp_2_41_10;
  wire pp_2_41_11;
  wire pp_2_42_0;
  wire pp_2_42_1;
  wire pp_2_42_2;
  wire pp_2_42_3;
  wire pp_2_42_4;
  wire pp_2_42_5;
  wire pp_2_42_6;
  wire pp_2_42_7;
  wire pp_2_42_8;
  wire pp_2_42_9;
  wire pp_2_43_0;
  wire pp_2_43_1;
  wire pp_2_43_2;
  wire pp_2_43_3;
  wire pp_2_43_4;
  wire pp_2_43_5;
  wire pp_2_43_6;
  wire pp_2_43_7;
  wire pp_2_43_8;
  wire pp_2_44_0;
  wire pp_2_44_1;
  wire pp_2_44_2;
  wire pp_2_44_3;
  wire pp_2_44_4;
  wire pp_2_44_5;
  wire pp_2_44_6;
  wire pp_2_44_7;
  wire pp_2_44_8;
  wire pp_2_44_9;
  wire pp_2_44_10;
  wire pp_2_44_11;
  wire pp_2_44_12;
  wire pp_2_44_13;
  wire pp_2_44_14;
  wire pp_2_44_15;
  wire pp_2_45_0;
  wire pp_2_45_1;
  wire pp_2_45_2;
  wire pp_2_45_3;
  wire pp_2_45_4;
  wire pp_2_45_5;
  wire pp_2_45_6;
  wire pp_2_45_7;
  wire pp_2_45_8;
  wire pp_2_46_0;
  wire pp_2_46_1;
  wire pp_2_46_2;
  wire pp_2_46_3;
  wire pp_2_46_4;
  wire pp_2_46_5;
  wire pp_2_46_6;
  wire pp_2_47_0;
  wire pp_2_47_1;
  wire pp_2_47_2;
  wire pp_2_47_3;
  wire pp_2_47_4;
  wire pp_2_47_5;
  wire pp_2_47_6;
  wire pp_2_47_7;
  wire pp_2_47_8;
  wire pp_2_48_0;
  wire pp_2_48_1;
  wire pp_2_48_2;
  wire pp_2_48_3;
  wire pp_2_48_4;
  wire pp_2_48_5;
  wire pp_2_48_6;
  wire pp_2_49_0;
  wire pp_2_49_1;
  wire pp_2_49_2;
  wire pp_2_49_3;
  wire pp_2_49_4;
  wire pp_2_49_5;
  wire pp_2_49_6;
  wire pp_2_49_7;
  wire pp_2_50_0;
  wire pp_2_50_1;
  wire pp_2_50_2;
  wire pp_2_50_3;
  wire pp_2_50_4;
  wire pp_2_50_5;
  wire pp_2_51_0;
  wire pp_2_51_1;
  wire pp_2_51_2;
  wire pp_2_51_3;
  wire pp_2_51_4;
  wire pp_2_51_5;
  wire pp_2_51_6;
  wire pp_2_52_0;
  wire pp_2_52_1;
  wire pp_2_52_2;
  wire pp_2_52_3;
  wire pp_2_52_4;
  wire pp_2_53_0;
  wire pp_2_53_1;
  wire pp_2_53_2;
  wire pp_2_53_3;
  wire pp_2_53_4;
  wire pp_2_53_5;
  wire pp_2_54_0;
  wire pp_2_54_1;
  wire pp_2_54_2;
  wire pp_2_54_3;
  wire pp_2_55_0;
  wire pp_2_55_1;
  wire pp_2_55_2;
  wire pp_2_55_3;
  wire pp_2_55_4;
  wire pp_2_56_0;
  wire pp_2_56_1;
  wire pp_2_56_2;
  wire pp_2_56_3;
  wire pp_2_56_4;
  wire pp_2_57_0;
  wire pp_2_57_1;
  wire pp_2_57_2;
  wire pp_2_57_3;
  wire pp_2_57_4;
  wire pp_2_58_0;
  wire pp_2_58_1;
  wire pp_2_58_2;
  wire pp_2_59_0;
  wire pp_2_59_1;
  wire pp_2_59_2;
  wire pp_2_59_3;
  wire pp_2_59_4;
  wire pp_2_59_5;
  wire pp_2_60_0;
  wire pp_2_61_0;
  wire pp_2_61_1;
  wire pp_2_61_2;
  wire pp_2_62_0;
  wire pp_3_0_0;
  wire pp_3_1_0;
  wire pp_3_1_1;
  wire pp_3_2_0;
  wire pp_3_2_1;
  wire pp_3_2_2;
  wire pp_3_3_0;
  wire pp_3_3_1;
  wire pp_3_3_2;
  wire pp_3_4_0;
  wire pp_3_4_1;
  wire pp_3_5_0;
  wire pp_3_5_1;
  wire pp_3_6_0;
  wire pp_3_6_1;
  wire pp_3_6_2;
  wire pp_3_6_3;
  wire pp_3_7_0;
  wire pp_3_7_1;
  wire pp_3_7_2;
  wire pp_3_7_3;
  wire pp_3_8_0;
  wire pp_3_8_1;
  wire pp_3_8_2;
  wire pp_3_8_3;
  wire pp_3_8_4;
  wire pp_3_8_5;
  wire pp_3_9_0;
  wire pp_3_9_1;
  wire pp_3_9_2;
  wire pp_3_10_0;
  wire pp_3_10_1;
  wire pp_3_10_2;
  wire pp_3_10_3;
  wire pp_3_10_4;
  wire pp_3_11_0;
  wire pp_3_11_1;
  wire pp_3_11_2;
  wire pp_3_11_3;
  wire pp_3_11_4;
  wire pp_3_11_5;
  wire pp_3_12_0;
  wire pp_3_12_1;
  wire pp_3_12_2;
  wire pp_3_13_0;
  wire pp_3_13_1;
  wire pp_3_13_2;
  wire pp_3_14_0;
  wire pp_3_14_1;
  wire pp_3_14_2;
  wire pp_3_14_3;
  wire pp_3_14_4;
  wire pp_3_14_5;
  wire pp_3_14_6;
  wire pp_3_14_7;
  wire pp_3_14_8;
  wire pp_3_15_0;
  wire pp_3_15_1;
  wire pp_3_15_2;
  wire pp_3_15_3;
  wire pp_3_15_4;
  wire pp_3_16_0;
  wire pp_3_16_1;
  wire pp_3_16_2;
  wire pp_3_16_3;
  wire pp_3_16_4;
  wire pp_3_16_5;
  wire pp_3_16_6;
  wire pp_3_16_7;
  wire pp_3_16_8;
  wire pp_3_17_0;
  wire pp_3_17_1;
  wire pp_3_17_2;
  wire pp_3_18_0;
  wire pp_3_18_1;
  wire pp_3_18_2;
  wire pp_3_18_3;
  wire pp_3_18_4;
  wire pp_3_18_5;
  wire pp_3_18_6;
  wire pp_3_18_7;
  wire pp_3_18_8;
  wire pp_3_18_9;
  wire pp_3_18_10;
  wire pp_3_19_0;
  wire pp_3_19_1;
  wire pp_3_19_2;
  wire pp_3_20_0;
  wire pp_3_20_1;
  wire pp_3_20_2;
  wire pp_3_20_3;
  wire pp_3_20_4;
  wire pp_3_20_5;
  wire pp_3_21_0;
  wire pp_3_21_1;
  wire pp_3_21_2;
  wire pp_3_21_3;
  wire pp_3_21_4;
  wire pp_3_21_5;
  wire pp_3_21_6;
  wire pp_3_21_7;
  wire pp_3_21_8;
  wire pp_3_22_0;
  wire pp_3_22_1;
  wire pp_3_22_2;
  wire pp_3_22_3;
  wire pp_3_22_4;
  wire pp_3_22_5;
  wire pp_3_22_6;
  wire pp_3_22_7;
  wire pp_3_22_8;
  wire pp_3_22_9;
  wire pp_3_22_10;
  wire pp_3_23_0;
  wire pp_3_23_1;
  wire pp_3_23_2;
  wire pp_3_23_3;
  wire pp_3_23_4;
  wire pp_3_23_5;
  wire pp_3_23_6;
  wire pp_3_23_7;
  wire pp_3_23_8;
  wire pp_3_24_0;
  wire pp_3_24_1;
  wire pp_3_24_2;
  wire pp_3_24_3;
  wire pp_3_24_4;
  wire pp_3_25_0;
  wire pp_3_25_1;
  wire pp_3_25_2;
  wire pp_3_25_3;
  wire pp_3_25_4;
  wire pp_3_25_5;
  wire pp_3_25_6;
  wire pp_3_25_7;
  wire pp_3_25_8;
  wire pp_3_25_9;
  wire pp_3_25_10;
  wire pp_3_25_11;
  wire pp_3_25_12;
  wire pp_3_25_13;
  wire pp_3_25_14;
  wire pp_3_26_0;
  wire pp_3_26_1;
  wire pp_3_26_2;
  wire pp_3_26_3;
  wire pp_3_26_4;
  wire pp_3_26_5;
  wire pp_3_26_6;
  wire pp_3_26_7;
  wire pp_3_27_0;
  wire pp_3_27_1;
  wire pp_3_27_2;
  wire pp_3_27_3;
  wire pp_3_27_4;
  wire pp_3_27_5;
  wire pp_3_27_6;
  wire pp_3_27_7;
  wire pp_3_27_8;
  wire pp_3_28_0;
  wire pp_3_28_1;
  wire pp_3_28_2;
  wire pp_3_28_3;
  wire pp_3_28_4;
  wire pp_3_28_5;
  wire pp_3_28_6;
  wire pp_3_28_7;
  wire pp_3_28_8;
  wire pp_3_29_0;
  wire pp_3_29_1;
  wire pp_3_29_2;
  wire pp_3_29_3;
  wire pp_3_29_4;
  wire pp_3_29_5;
  wire pp_3_29_6;
  wire pp_3_29_7;
  wire pp_3_29_8;
  wire pp_3_30_0;
  wire pp_3_30_1;
  wire pp_3_30_2;
  wire pp_3_30_3;
  wire pp_3_30_4;
  wire pp_3_30_5;
  wire pp_3_30_6;
  wire pp_3_30_7;
  wire pp_3_30_8;
  wire pp_3_31_0;
  wire pp_3_31_1;
  wire pp_3_31_2;
  wire pp_3_31_3;
  wire pp_3_31_4;
  wire pp_3_31_5;
  wire pp_3_31_6;
  wire pp_3_31_7;
  wire pp_3_31_8;
  wire pp_3_32_0;
  wire pp_3_32_1;
  wire pp_3_32_2;
  wire pp_3_32_3;
  wire pp_3_32_4;
  wire pp_3_32_5;
  wire pp_3_32_6;
  wire pp_3_32_7;
  wire pp_3_32_8;
  wire pp_3_32_9;
  wire pp_3_32_10;
  wire pp_3_33_0;
  wire pp_3_33_1;
  wire pp_3_33_2;
  wire pp_3_33_3;
  wire pp_3_33_4;
  wire pp_3_33_5;
  wire pp_3_33_6;
  wire pp_3_33_7;
  wire pp_3_33_8;
  wire pp_3_34_0;
  wire pp_3_34_1;
  wire pp_3_34_2;
  wire pp_3_34_3;
  wire pp_3_34_4;
  wire pp_3_34_5;
  wire pp_3_34_6;
  wire pp_3_34_7;
  wire pp_3_34_8;
  wire pp_3_34_9;
  wire pp_3_35_0;
  wire pp_3_35_1;
  wire pp_3_35_2;
  wire pp_3_35_3;
  wire pp_3_35_4;
  wire pp_3_35_5;
  wire pp_3_35_6;
  wire pp_3_35_7;
  wire pp_3_35_8;
  wire pp_3_35_9;
  wire pp_3_36_0;
  wire pp_3_36_1;
  wire pp_3_36_2;
  wire pp_3_36_3;
  wire pp_3_36_4;
  wire pp_3_36_5;
  wire pp_3_36_6;
  wire pp_3_36_7;
  wire pp_3_37_0;
  wire pp_3_37_1;
  wire pp_3_37_2;
  wire pp_3_37_3;
  wire pp_3_37_4;
  wire pp_3_37_5;
  wire pp_3_37_6;
  wire pp_3_37_7;
  wire pp_3_37_8;
  wire pp_3_38_0;
  wire pp_3_38_1;
  wire pp_3_38_2;
  wire pp_3_38_3;
  wire pp_3_38_4;
  wire pp_3_38_5;
  wire pp_3_38_6;
  wire pp_3_38_7;
  wire pp_3_38_8;
  wire pp_3_39_0;
  wire pp_3_39_1;
  wire pp_3_39_2;
  wire pp_3_39_3;
  wire pp_3_39_4;
  wire pp_3_39_5;
  wire pp_3_39_6;
  wire pp_3_39_7;
  wire pp_3_39_8;
  wire pp_3_40_0;
  wire pp_3_40_1;
  wire pp_3_40_2;
  wire pp_3_40_3;
  wire pp_3_40_4;
  wire pp_3_40_5;
  wire pp_3_40_6;
  wire pp_3_41_0;
  wire pp_3_41_1;
  wire pp_3_41_2;
  wire pp_3_41_3;
  wire pp_3_41_4;
  wire pp_3_41_5;
  wire pp_3_41_6;
  wire pp_3_41_7;
  wire pp_3_41_8;
  wire pp_3_41_9;
  wire pp_3_41_10;
  wire pp_3_41_11;
  wire pp_3_42_0;
  wire pp_3_42_1;
  wire pp_3_42_2;
  wire pp_3_42_3;
  wire pp_3_42_4;
  wire pp_3_42_5;
  wire pp_3_43_0;
  wire pp_3_43_1;
  wire pp_3_43_2;
  wire pp_3_43_3;
  wire pp_3_43_4;
  wire pp_3_43_5;
  wire pp_3_44_0;
  wire pp_3_44_1;
  wire pp_3_44_2;
  wire pp_3_44_3;
  wire pp_3_44_4;
  wire pp_3_44_5;
  wire pp_3_44_6;
  wire pp_3_44_7;
  wire pp_3_44_8;
  wire pp_3_45_0;
  wire pp_3_45_1;
  wire pp_3_45_2;
  wire pp_3_45_3;
  wire pp_3_45_4;
  wire pp_3_45_5;
  wire pp_3_45_6;
  wire pp_3_45_7;
  wire pp_3_45_8;
  wire pp_3_45_9;
  wire pp_3_46_0;
  wire pp_3_46_1;
  wire pp_3_46_2;
  wire pp_3_46_3;
  wire pp_3_46_4;
  wire pp_3_46_5;
  wire pp_3_46_6;
  wire pp_3_46_7;
  wire pp_3_46_8;
  wire pp_3_47_0;
  wire pp_3_47_1;
  wire pp_3_47_2;
  wire pp_3_48_0;
  wire pp_3_48_1;
  wire pp_3_48_2;
  wire pp_3_48_3;
  wire pp_3_48_4;
  wire pp_3_48_5;
  wire pp_3_49_0;
  wire pp_3_49_1;
  wire pp_3_49_2;
  wire pp_3_49_3;
  wire pp_3_49_4;
  wire pp_3_49_5;
  wire pp_3_50_0;
  wire pp_3_50_1;
  wire pp_3_50_2;
  wire pp_3_50_3;
  wire pp_3_50_4;
  wire pp_3_50_5;
  wire pp_3_51_0;
  wire pp_3_51_1;
  wire pp_3_51_2;
  wire pp_3_51_3;
  wire pp_3_51_4;
  wire pp_3_51_5;
  wire pp_3_52_0;
  wire pp_3_52_1;
  wire pp_3_52_2;
  wire pp_3_52_3;
  wire pp_3_53_0;
  wire pp_3_53_1;
  wire pp_3_53_2;
  wire pp_3_54_0;
  wire pp_3_54_1;
  wire pp_3_54_2;
  wire pp_3_54_3;
  wire pp_3_54_4;
  wire pp_3_54_5;
  wire pp_3_55_0;
  wire pp_3_55_1;
  wire pp_3_55_2;
  wire pp_3_56_0;
  wire pp_3_56_1;
  wire pp_3_56_2;
  wire pp_3_56_3;
  wire pp_3_56_4;
  wire pp_3_56_5;
  wire pp_3_57_0;
  wire pp_3_57_1;
  wire pp_3_57_2;
  wire pp_3_58_0;
  wire pp_3_58_1;
  wire pp_3_59_0;
  wire pp_3_59_1;
  wire pp_3_59_2;
  wire pp_3_60_0;
  wire pp_3_60_1;
  wire pp_3_60_2;
  wire pp_3_61_0;
  wire pp_3_62_0;
  wire pp_3_62_1;
  wire pp_4_0_0;
  wire pp_4_1_0;
  wire pp_4_1_1;
  wire pp_4_2_0;
  wire pp_4_2_1;
  wire pp_4_2_2;
  wire pp_4_3_0;
  wire pp_4_4_0;
  wire pp_4_4_1;
  wire pp_4_5_0;
  wire pp_4_5_1;
  wire pp_4_6_0;
  wire pp_4_6_1;
  wire pp_4_6_2;
  wire pp_4_7_0;
  wire pp_4_7_1;
  wire pp_4_7_2;
  wire pp_4_8_0;
  wire pp_4_8_1;
  wire pp_4_8_2;
  wire pp_4_9_0;
  wire pp_4_9_1;
  wire pp_4_9_2;
  wire pp_4_10_0;
  wire pp_4_10_1;
  wire pp_4_10_2;
  wire pp_4_11_0;
  wire pp_4_11_1;
  wire pp_4_11_2;
  wire pp_4_11_3;
  wire pp_4_12_0;
  wire pp_4_12_1;
  wire pp_4_12_2;
  wire pp_4_13_0;
  wire pp_4_13_1;
  wire pp_4_14_0;
  wire pp_4_14_1;
  wire pp_4_14_2;
  wire pp_4_14_3;
  wire pp_4_15_0;
  wire pp_4_15_1;
  wire pp_4_15_2;
  wire pp_4_15_3;
  wire pp_4_15_4;
  wire pp_4_15_5;
  wire pp_4_16_0;
  wire pp_4_16_1;
  wire pp_4_16_2;
  wire pp_4_16_3;
  wire pp_4_17_0;
  wire pp_4_17_1;
  wire pp_4_17_2;
  wire pp_4_17_3;
  wire pp_4_18_0;
  wire pp_4_18_1;
  wire pp_4_18_2;
  wire pp_4_18_3;
  wire pp_4_18_4;
  wire pp_4_18_5;
  wire pp_4_19_0;
  wire pp_4_19_1;
  wire pp_4_19_2;
  wire pp_4_19_3;
  wire pp_4_20_0;
  wire pp_4_20_1;
  wire pp_4_20_2;
  wire pp_4_21_0;
  wire pp_4_21_1;
  wire pp_4_21_2;
  wire pp_4_21_3;
  wire pp_4_21_4;
  wire pp_4_22_0;
  wire pp_4_22_1;
  wire pp_4_22_2;
  wire pp_4_22_3;
  wire pp_4_22_4;
  wire pp_4_22_5;
  wire pp_4_22_6;
  wire pp_4_22_7;
  wire pp_4_23_0;
  wire pp_4_23_1;
  wire pp_4_23_2;
  wire pp_4_23_3;
  wire pp_4_23_4;
  wire pp_4_23_5;
  wire pp_4_24_0;
  wire pp_4_24_1;
  wire pp_4_24_2;
  wire pp_4_24_3;
  wire pp_4_24_4;
  wire pp_4_24_5;
  wire pp_4_25_0;
  wire pp_4_25_1;
  wire pp_4_25_2;
  wire pp_4_25_3;
  wire pp_4_25_4;
  wire pp_4_25_5;
  wire pp_4_26_0;
  wire pp_4_26_1;
  wire pp_4_26_2;
  wire pp_4_26_3;
  wire pp_4_26_4;
  wire pp_4_26_5;
  wire pp_4_26_6;
  wire pp_4_26_7;
  wire pp_4_26_8;
  wire pp_4_27_0;
  wire pp_4_27_1;
  wire pp_4_27_2;
  wire pp_4_27_3;
  wire pp_4_27_4;
  wire pp_4_28_0;
  wire pp_4_28_1;
  wire pp_4_28_2;
  wire pp_4_28_3;
  wire pp_4_28_4;
  wire pp_4_28_5;
  wire pp_4_29_0;
  wire pp_4_29_1;
  wire pp_4_29_2;
  wire pp_4_29_3;
  wire pp_4_29_4;
  wire pp_4_29_5;
  wire pp_4_30_0;
  wire pp_4_30_1;
  wire pp_4_30_2;
  wire pp_4_30_3;
  wire pp_4_30_4;
  wire pp_4_30_5;
  wire pp_4_31_0;
  wire pp_4_31_1;
  wire pp_4_31_2;
  wire pp_4_31_3;
  wire pp_4_31_4;
  wire pp_4_31_5;
  wire pp_4_32_0;
  wire pp_4_32_1;
  wire pp_4_32_2;
  wire pp_4_32_3;
  wire pp_4_32_4;
  wire pp_4_32_5;
  wire pp_4_32_6;
  wire pp_4_32_7;
  wire pp_4_33_0;
  wire pp_4_33_1;
  wire pp_4_33_2;
  wire pp_4_33_3;
  wire pp_4_33_4;
  wire pp_4_33_5;
  wire pp_4_34_0;
  wire pp_4_34_1;
  wire pp_4_34_2;
  wire pp_4_34_3;
  wire pp_4_34_4;
  wire pp_4_34_5;
  wire pp_4_34_6;
  wire pp_4_35_0;
  wire pp_4_35_1;
  wire pp_4_35_2;
  wire pp_4_35_3;
  wire pp_4_35_4;
  wire pp_4_35_5;
  wire pp_4_35_6;
  wire pp_4_35_7;
  wire pp_4_35_8;
  wire pp_4_36_0;
  wire pp_4_36_1;
  wire pp_4_36_2;
  wire pp_4_36_3;
  wire pp_4_36_4;
  wire pp_4_36_5;
  wire pp_4_37_0;
  wire pp_4_37_1;
  wire pp_4_37_2;
  wire pp_4_37_3;
  wire pp_4_37_4;
  wire pp_4_37_5;
  wire pp_4_37_6;
  wire pp_4_37_7;
  wire pp_4_37_8;
  wire pp_4_38_0;
  wire pp_4_38_1;
  wire pp_4_38_2;
  wire pp_4_38_3;
  wire pp_4_38_4;
  wire pp_4_38_5;
  wire pp_4_39_0;
  wire pp_4_39_1;
  wire pp_4_39_2;
  wire pp_4_39_3;
  wire pp_4_39_4;
  wire pp_4_40_0;
  wire pp_4_40_1;
  wire pp_4_40_2;
  wire pp_4_40_3;
  wire pp_4_40_4;
  wire pp_4_40_5;
  wire pp_4_41_0;
  wire pp_4_41_1;
  wire pp_4_41_2;
  wire pp_4_41_3;
  wire pp_4_41_4;
  wire pp_4_41_5;
  wire pp_4_42_0;
  wire pp_4_42_1;
  wire pp_4_42_2;
  wire pp_4_42_3;
  wire pp_4_42_4;
  wire pp_4_42_5;
  wire pp_4_42_6;
  wire pp_4_42_7;
  wire pp_4_43_0;
  wire pp_4_43_1;
  wire pp_4_43_2;
  wire pp_4_44_0;
  wire pp_4_44_1;
  wire pp_4_44_2;
  wire pp_4_44_3;
  wire pp_4_44_4;
  wire pp_4_45_0;
  wire pp_4_45_1;
  wire pp_4_45_2;
  wire pp_4_45_3;
  wire pp_4_45_4;
  wire pp_4_45_5;
  wire pp_4_45_6;
  wire pp_4_46_0;
  wire pp_4_46_1;
  wire pp_4_46_2;
  wire pp_4_46_3;
  wire pp_4_46_4;
  wire pp_4_46_5;
  wire pp_4_46_6;
  wire pp_4_46_7;
  wire pp_4_47_0;
  wire pp_4_47_1;
  wire pp_4_47_2;
  wire pp_4_48_0;
  wire pp_4_48_1;
  wire pp_4_48_2;
  wire pp_4_49_0;
  wire pp_4_49_1;
  wire pp_4_49_2;
  wire pp_4_49_3;
  wire pp_4_50_0;
  wire pp_4_50_1;
  wire pp_4_50_2;
  wire pp_4_50_3;
  wire pp_4_50_4;
  wire pp_4_50_5;
  wire pp_4_51_0;
  wire pp_4_51_1;
  wire pp_4_51_2;
  wire pp_4_52_0;
  wire pp_4_52_1;
  wire pp_4_52_2;
  wire pp_4_52_3;
  wire pp_4_52_4;
  wire pp_4_52_5;
  wire pp_4_53_0;
  wire pp_4_54_0;
  wire pp_4_54_1;
  wire pp_4_54_2;
  wire pp_4_55_0;
  wire pp_4_55_1;
  wire pp_4_55_2;
  wire pp_4_56_0;
  wire pp_4_56_1;
  wire pp_4_56_2;
  wire pp_4_57_0;
  wire pp_4_57_1;
  wire pp_4_57_2;
  wire pp_4_58_0;
  wire pp_4_58_1;
  wire pp_4_58_2;
  wire pp_4_59_0;
  wire pp_4_60_0;
  wire pp_4_60_1;
  wire pp_4_61_0;
  wire pp_4_61_1;
  wire pp_4_62_0;
  wire pp_4_62_1;
  wire pp_5_0_0;
  wire pp_5_1_0;
  wire pp_5_1_1;
  wire pp_5_2_0;
  wire pp_5_2_1;
  wire pp_5_3_0;
  wire pp_5_3_1;
  wire pp_5_4_0;
  wire pp_5_4_1;
  wire pp_5_5_0;
  wire pp_5_5_1;
  wire pp_5_6_0;
  wire pp_5_6_1;
  wire pp_5_6_2;
  wire pp_5_7_0;
  wire pp_5_8_0;
  wire pp_5_8_1;
  wire pp_5_9_0;
  wire pp_5_9_1;
  wire pp_5_10_0;
  wire pp_5_10_1;
  wire pp_5_11_0;
  wire pp_5_11_1;
  wire pp_5_11_2;
  wire pp_5_11_3;
  wire pp_5_12_0;
  wire pp_5_12_1;
  wire pp_5_13_0;
  wire pp_5_13_1;
  wire pp_5_13_2;
  wire pp_5_14_0;
  wire pp_5_14_1;
  wire pp_5_15_0;
  wire pp_5_15_1;
  wire pp_5_15_2;
  wire pp_5_16_0;
  wire pp_5_16_1;
  wire pp_5_16_2;
  wire pp_5_16_3;
  wire pp_5_16_4;
  wire pp_5_16_5;
  wire pp_5_17_0;
  wire pp_5_17_1;
  wire pp_5_18_0;
  wire pp_5_18_1;
  wire pp_5_18_2;
  wire pp_5_19_0;
  wire pp_5_19_1;
  wire pp_5_19_2;
  wire pp_5_19_3;
  wire pp_5_19_4;
  wire pp_5_19_5;
  wire pp_5_20_0;
  wire pp_5_21_0;
  wire pp_5_21_1;
  wire pp_5_21_2;
  wire pp_5_22_0;
  wire pp_5_22_1;
  wire pp_5_22_2;
  wire pp_5_22_3;
  wire pp_5_22_4;
  wire pp_5_22_5;
  wire pp_5_23_0;
  wire pp_5_23_1;
  wire pp_5_23_2;
  wire pp_5_23_3;
  wire pp_5_24_0;
  wire pp_5_24_1;
  wire pp_5_24_2;
  wire pp_5_24_3;
  wire pp_5_25_0;
  wire pp_5_25_1;
  wire pp_5_25_2;
  wire pp_5_25_3;
  wire pp_5_26_0;
  wire pp_5_26_1;
  wire pp_5_26_2;
  wire pp_5_26_3;
  wire pp_5_26_4;
  wire pp_5_26_5;
  wire pp_5_26_6;
  wire pp_5_26_7;
  wire pp_5_26_8;
  wire pp_5_27_0;
  wire pp_5_27_1;
  wire pp_5_27_2;
  wire pp_5_27_3;
  wire pp_5_28_0;
  wire pp_5_28_1;
  wire pp_5_28_2;
  wire pp_5_29_0;
  wire pp_5_29_1;
  wire pp_5_29_2;
  wire pp_5_29_3;
  wire pp_5_29_4;
  wire pp_5_30_0;
  wire pp_5_30_1;
  wire pp_5_30_2;
  wire pp_5_30_3;
  wire pp_5_31_0;
  wire pp_5_31_1;
  wire pp_5_31_2;
  wire pp_5_31_3;
  wire pp_5_31_4;
  wire pp_5_31_5;
  wire pp_5_32_0;
  wire pp_5_32_1;
  wire pp_5_32_2;
  wire pp_5_32_3;
  wire pp_5_32_4;
  wire pp_5_33_0;
  wire pp_5_33_1;
  wire pp_5_33_2;
  wire pp_5_33_3;
  wire pp_5_34_0;
  wire pp_5_34_1;
  wire pp_5_34_2;
  wire pp_5_34_3;
  wire pp_5_34_4;
  wire pp_5_34_5;
  wire pp_5_34_6;
  wire pp_5_34_7;
  wire pp_5_34_8;
  wire pp_5_35_0;
  wire pp_5_35_1;
  wire pp_5_35_2;
  wire pp_5_36_0;
  wire pp_5_36_1;
  wire pp_5_36_2;
  wire pp_5_36_3;
  wire pp_5_36_4;
  wire pp_5_36_5;
  wire pp_5_36_6;
  wire pp_5_36_7;
  wire pp_5_36_8;
  wire pp_5_37_0;
  wire pp_5_37_1;
  wire pp_5_37_2;
  wire pp_5_38_0;
  wire pp_5_38_1;
  wire pp_5_38_2;
  wire pp_5_38_3;
  wire pp_5_38_4;
  wire pp_5_38_5;
  wire pp_5_38_6;
  wire pp_5_38_7;
  wire pp_5_38_8;
  wire pp_5_39_0;
  wire pp_5_39_1;
  wire pp_5_39_2;
  wire pp_5_40_0;
  wire pp_5_40_1;
  wire pp_5_40_2;
  wire pp_5_41_0;
  wire pp_5_41_1;
  wire pp_5_41_2;
  wire pp_5_41_3;
  wire pp_5_41_4;
  wire pp_5_41_5;
  wire pp_5_41_6;
  wire pp_5_41_7;
  wire pp_5_42_0;
  wire pp_5_42_1;
  wire pp_5_42_2;
  wire pp_5_42_3;
  wire pp_5_43_0;
  wire pp_5_43_1;
  wire pp_5_43_2;
  wire pp_5_44_0;
  wire pp_5_44_1;
  wire pp_5_44_2;
  wire pp_5_44_3;
  wire pp_5_44_4;
  wire pp_5_44_5;
  wire pp_5_45_0;
  wire pp_5_45_1;
  wire pp_5_45_2;
  wire pp_5_46_0;
  wire pp_5_46_1;
  wire pp_5_46_2;
  wire pp_5_46_3;
  wire pp_5_46_4;
  wire pp_5_46_5;
  wire pp_5_47_0;
  wire pp_5_47_1;
  wire pp_5_47_2;
  wire pp_5_48_0;
  wire pp_5_48_1;
  wire pp_5_48_2;
  wire pp_5_48_3;
  wire pp_5_49_0;
  wire pp_5_49_1;
  wire pp_5_50_0;
  wire pp_5_50_1;
  wire pp_5_50_2;
  wire pp_5_50_3;
  wire pp_5_50_4;
  wire pp_5_50_5;
  wire pp_5_50_6;
  wire pp_5_51_0;
  wire pp_5_52_0;
  wire pp_5_52_1;
  wire pp_5_52_2;
  wire pp_5_52_3;
  wire pp_5_52_4;
  wire pp_5_52_5;
  wire pp_5_52_6;
  wire pp_5_53_0;
  wire pp_5_54_0;
  wire pp_5_54_1;
  wire pp_5_54_2;
  wire pp_5_55_0;
  wire pp_5_55_1;
  wire pp_5_55_2;
  wire pp_5_56_0;
  wire pp_5_56_1;
  wire pp_5_56_2;
  wire pp_5_57_0;
  wire pp_5_58_0;
  wire pp_5_58_1;
  wire pp_5_59_0;
  wire pp_5_59_1;
  wire pp_5_60_0;
  wire pp_5_60_1;
  wire pp_5_61_0;
  wire pp_5_61_1;
  wire pp_5_62_0;
  wire pp_5_62_1;
  wire pp_6_0_0;
  wire pp_6_1_0;
  wire pp_6_1_1;
  wire pp_6_2_0;
  wire pp_6_2_1;
  wire pp_6_3_0;
  wire pp_6_3_1;
  wire pp_6_4_0;
  wire pp_6_4_1;
  wire pp_6_5_0;
  wire pp_6_5_1;
  wire pp_6_6_0;
  wire pp_6_6_1;
  wire pp_6_6_2;
  wire pp_6_7_0;
  wire pp_6_8_0;
  wire pp_6_8_1;
  wire pp_6_9_0;
  wire pp_6_9_1;
  wire pp_6_10_0;
  wire pp_6_10_1;
  wire pp_6_11_0;
  wire pp_6_11_1;
  wire pp_6_11_2;
  wire pp_6_11_3;
  wire pp_6_12_0;
  wire pp_6_13_0;
  wire pp_6_13_1;
  wire pp_6_14_0;
  wire pp_6_14_1;
  wire pp_6_14_2;
  wire pp_6_15_0;
  wire pp_6_16_0;
  wire pp_6_16_1;
  wire pp_6_16_2;
  wire pp_6_17_0;
  wire pp_6_17_1;
  wire pp_6_17_2;
  wire pp_6_18_0;
  wire pp_6_18_1;
  wire pp_6_19_0;
  wire pp_6_19_1;
  wire pp_6_19_2;
  wire pp_6_20_0;
  wire pp_6_20_1;
  wire pp_6_20_2;
  wire pp_6_21_0;
  wire pp_6_21_1;
  wire pp_6_21_2;
  wire pp_6_22_0;
  wire pp_6_22_1;
  wire pp_6_23_0;
  wire pp_6_23_1;
  wire pp_6_23_2;
  wire pp_6_23_3;
  wire pp_6_24_0;
  wire pp_6_24_1;
  wire pp_6_24_2;
  wire pp_6_25_0;
  wire pp_6_25_1;
  wire pp_6_25_2;
  wire pp_6_25_3;
  wire pp_6_26_0;
  wire pp_6_26_1;
  wire pp_6_26_2;
  wire pp_6_26_3;
  wire pp_6_27_0;
  wire pp_6_27_1;
  wire pp_6_27_2;
  wire pp_6_27_3;
  wire pp_6_27_4;
  wire pp_6_28_0;
  wire pp_6_28_1;
  wire pp_6_29_0;
  wire pp_6_29_1;
  wire pp_6_29_2;
  wire pp_6_29_3;
  wire pp_6_30_0;
  wire pp_6_30_1;
  wire pp_6_30_2;
  wire pp_6_31_0;
  wire pp_6_31_1;
  wire pp_6_31_2;
  wire pp_6_32_0;
  wire pp_6_32_1;
  wire pp_6_32_2;
  wire pp_6_32_3;
  wire pp_6_32_4;
  wire pp_6_33_0;
  wire pp_6_33_1;
  wire pp_6_33_2;
  wire pp_6_34_0;
  wire pp_6_34_1;
  wire pp_6_34_2;
  wire pp_6_34_3;
  wire pp_6_35_0;
  wire pp_6_35_1;
  wire pp_6_35_2;
  wire pp_6_35_3;
  wire pp_6_36_0;
  wire pp_6_36_1;
  wire pp_6_36_2;
  wire pp_6_36_3;
  wire pp_6_37_0;
  wire pp_6_37_1;
  wire pp_6_37_2;
  wire pp_6_37_3;
  wire pp_6_38_0;
  wire pp_6_38_1;
  wire pp_6_38_2;
  wire pp_6_38_3;
  wire pp_6_39_0;
  wire pp_6_39_1;
  wire pp_6_39_2;
  wire pp_6_39_3;
  wire pp_6_40_0;
  wire pp_6_40_1;
  wire pp_6_41_0;
  wire pp_6_41_1;
  wire pp_6_41_2;
  wire pp_6_41_3;
  wire pp_6_41_4;
  wire pp_6_41_5;
  wire pp_6_41_6;
  wire pp_6_42_0;
  wire pp_6_42_1;
  wire pp_6_42_2;
  wire pp_6_43_0;
  wire pp_6_43_1;
  wire pp_6_44_0;
  wire pp_6_44_1;
  wire pp_6_44_2;
  wire pp_6_45_0;
  wire pp_6_45_1;
  wire pp_6_45_2;
  wire pp_6_45_3;
  wire pp_6_45_4;
  wire pp_6_46_0;
  wire pp_6_46_1;
  wire pp_6_47_0;
  wire pp_6_47_1;
  wire pp_6_47_2;
  wire pp_6_48_0;
  wire pp_6_48_1;
  wire pp_6_48_2;
  wire pp_6_49_0;
  wire pp_6_49_1;
  wire pp_6_49_2;
  wire pp_6_50_0;
  wire pp_6_50_1;
  wire pp_6_50_2;
  wire pp_6_51_0;
  wire pp_6_51_1;
  wire pp_6_51_2;
  wire pp_6_52_0;
  wire pp_6_52_1;
  wire pp_6_52_2;
  wire pp_6_53_0;
  wire pp_6_53_1;
  wire pp_6_53_2;
  wire pp_6_54_0;
  wire pp_6_55_0;
  wire pp_6_55_1;
  wire pp_6_56_0;
  wire pp_6_56_1;
  wire pp_6_57_0;
  wire pp_6_57_1;
  wire pp_6_58_0;
  wire pp_6_58_1;
  wire pp_6_59_0;
  wire pp_6_59_1;
  wire pp_6_60_0;
  wire pp_6_60_1;
  wire pp_6_61_0;
  wire pp_6_61_1;
  wire pp_6_62_0;
  wire pp_6_62_1;
  wire pp_7_0_0;
  wire pp_7_1_0;
  wire pp_7_1_1;
  wire pp_7_2_0;
  wire pp_7_2_1;
  wire pp_7_3_0;
  wire pp_7_3_1;
  wire pp_7_4_0;
  wire pp_7_4_1;
  wire pp_7_5_0;
  wire pp_7_5_1;
  wire pp_7_6_0;
  wire pp_7_6_1;
  wire pp_7_6_2;
  wire pp_7_7_0;
  wire pp_7_8_0;
  wire pp_7_8_1;
  wire pp_7_9_0;
  wire pp_7_9_1;
  wire pp_7_10_0;
  wire pp_7_10_1;
  wire pp_7_11_0;
  wire pp_7_11_1;
  wire pp_7_12_0;
  wire pp_7_12_1;
  wire pp_7_13_0;
  wire pp_7_13_1;
  wire pp_7_14_0;
  wire pp_7_14_1;
  wire pp_7_15_0;
  wire pp_7_15_1;
  wire pp_7_16_0;
  wire pp_7_16_1;
  wire pp_7_17_0;
  wire pp_7_17_1;
  wire pp_7_17_2;
  wire pp_7_17_3;
  wire pp_7_18_0;
  wire pp_7_18_1;
  wire pp_7_19_0;
  wire pp_7_20_0;
  wire pp_7_20_1;
  wire pp_7_20_2;
  wire pp_7_20_3;
  wire pp_7_21_0;
  wire pp_7_21_1;
  wire pp_7_21_2;
  wire pp_7_22_0;
  wire pp_7_23_0;
  wire pp_7_23_1;
  wire pp_7_23_2;
  wire pp_7_24_0;
  wire pp_7_24_1;
  wire pp_7_25_0;
  wire pp_7_25_1;
  wire pp_7_25_2;
  wire pp_7_26_0;
  wire pp_7_26_1;
  wire pp_7_26_2;
  wire pp_7_27_0;
  wire pp_7_27_1;
  wire pp_7_27_2;
  wire pp_7_28_0;
  wire pp_7_28_1;
  wire pp_7_28_2;
  wire pp_7_29_0;
  wire pp_7_29_1;
  wire pp_7_29_2;
  wire pp_7_30_0;
  wire pp_7_30_1;
  wire pp_7_30_2;
  wire pp_7_31_0;
  wire pp_7_31_1;
  wire pp_7_31_2;
  wire pp_7_32_0;
  wire pp_7_32_1;
  wire pp_7_32_2;
  wire pp_7_33_0;
  wire pp_7_33_1;
  wire pp_7_33_2;
  wire pp_7_34_0;
  wire pp_7_34_1;
  wire pp_7_34_2;
  wire pp_7_35_0;
  wire pp_7_35_1;
  wire pp_7_35_2;
  wire pp_7_36_0;
  wire pp_7_36_1;
  wire pp_7_36_2;
  wire pp_7_37_0;
  wire pp_7_37_1;
  wire pp_7_37_2;
  wire pp_7_38_0;
  wire pp_7_38_1;
  wire pp_7_38_2;
  wire pp_7_39_0;
  wire pp_7_39_1;
  wire pp_7_39_2;
  wire pp_7_40_0;
  wire pp_7_40_1;
  wire pp_7_40_2;
  wire pp_7_41_0;
  wire pp_7_41_1;
  wire pp_7_41_2;
  wire pp_7_42_0;
  wire pp_7_42_1;
  wire pp_7_42_2;
  wire pp_7_43_0;
  wire pp_7_43_1;
  wire pp_7_43_2;
  wire pp_7_44_0;
  wire pp_7_45_0;
  wire pp_7_45_1;
  wire pp_7_45_2;
  wire pp_7_45_3;
  wire pp_7_46_0;
  wire pp_7_46_1;
  wire pp_7_46_2;
  wire pp_7_47_0;
  wire pp_7_48_0;
  wire pp_7_48_1;
  wire pp_7_49_0;
  wire pp_7_49_1;
  wire pp_7_49_2;
  wire pp_7_49_3;
  wire pp_7_50_0;
  wire pp_7_50_1;
  wire pp_7_50_2;
  wire pp_7_51_0;
  wire pp_7_52_0;
  wire pp_7_52_1;
  wire pp_7_53_0;
  wire pp_7_53_1;
  wire pp_7_53_2;
  wire pp_7_53_3;
  wire pp_7_54_0;
  wire pp_7_55_0;
  wire pp_7_55_1;
  wire pp_7_56_0;
  wire pp_7_56_1;
  wire pp_7_57_0;
  wire pp_7_57_1;
  wire pp_7_58_0;
  wire pp_7_58_1;
  wire pp_7_59_0;
  wire pp_7_59_1;
  wire pp_7_60_0;
  wire pp_7_60_1;
  wire pp_7_61_0;
  wire pp_7_61_1;
  wire pp_7_62_0;
  wire pp_7_62_1;
  wire pp_8_0_0;
  wire pp_8_1_0;
  wire pp_8_1_1;
  wire pp_8_2_0;
  wire pp_8_2_1;
  wire pp_8_3_0;
  wire pp_8_3_1;
  wire pp_8_4_0;
  wire pp_8_4_1;
  wire pp_8_5_0;
  wire pp_8_5_1;
  wire pp_8_6_0;
  wire pp_8_6_1;
  wire pp_8_7_0;
  wire pp_8_7_1;
  wire pp_8_8_0;
  wire pp_8_8_1;
  wire pp_8_9_0;
  wire pp_8_9_1;
  wire pp_8_10_0;
  wire pp_8_10_1;
  wire pp_8_11_0;
  wire pp_8_11_1;
  wire pp_8_12_0;
  wire pp_8_12_1;
  wire pp_8_13_0;
  wire pp_8_13_1;
  wire pp_8_14_0;
  wire pp_8_14_1;
  wire pp_8_15_0;
  wire pp_8_15_1;
  wire pp_8_16_0;
  wire pp_8_16_1;
  wire pp_8_17_0;
  wire pp_8_17_1;
  wire pp_8_18_0;
  wire pp_8_18_1;
  wire pp_8_19_0;
  wire pp_8_19_1;
  wire pp_8_20_0;
  wire pp_8_20_1;
  wire pp_8_21_0;
  wire pp_8_21_1;
  wire pp_8_22_0;
  wire pp_8_22_1;
  wire pp_8_23_0;
  wire pp_8_23_1;
  wire pp_8_24_0;
  wire pp_8_24_1;
  wire pp_8_25_0;
  wire pp_8_25_1;
  wire pp_8_26_0;
  wire pp_8_26_1;
  wire pp_8_27_0;
  wire pp_8_27_1;
  wire pp_8_28_0;
  wire pp_8_28_1;
  wire pp_8_29_0;
  wire pp_8_29_1;
  wire pp_8_30_0;
  wire pp_8_30_1;
  wire pp_8_31_0;
  wire pp_8_31_1;
  wire pp_8_32_0;
  wire pp_8_32_1;
  wire pp_8_33_0;
  wire pp_8_33_1;
  wire pp_8_34_0;
  wire pp_8_34_1;
  wire pp_8_35_0;
  wire pp_8_35_1;
  wire pp_8_36_0;
  wire pp_8_36_1;
  wire pp_8_37_0;
  wire pp_8_37_1;
  wire pp_8_38_0;
  wire pp_8_38_1;
  wire pp_8_39_0;
  wire pp_8_39_1;
  wire pp_8_40_0;
  wire pp_8_40_1;
  wire pp_8_41_0;
  wire pp_8_41_1;
  wire pp_8_42_0;
  wire pp_8_42_1;
  wire pp_8_43_0;
  wire pp_8_43_1;
  wire pp_8_44_0;
  wire pp_8_44_1;
  wire pp_8_45_0;
  wire pp_8_45_1;
  wire pp_8_46_0;
  wire pp_8_46_1;
  wire pp_8_47_0;
  wire pp_8_47_1;
  wire pp_8_48_0;
  wire pp_8_48_1;
  wire pp_8_49_0;
  wire pp_8_49_1;
  wire pp_8_50_0;
  wire pp_8_50_1;
  wire pp_8_51_0;
  wire pp_8_51_1;
  wire pp_8_52_0;
  wire pp_8_52_1;
  wire pp_8_53_0;
  wire pp_8_53_1;
  wire pp_8_54_0;
  wire pp_8_54_1;
  wire pp_8_55_0;
  wire pp_8_55_1;
  wire pp_8_56_0;
  wire pp_8_56_1;
  wire pp_8_57_0;
  wire pp_8_57_1;
  wire pp_8_58_0;
  wire pp_8_58_1;
  wire pp_8_59_0;
  wire pp_8_59_1;
  wire pp_8_60_0;
  wire pp_8_60_1;
  wire pp_8_61_0;
  wire pp_8_61_1;
  wire pp_8_62_0;
  wire pp_8_62_1;
  assign pp_0_0_0 = pp_0_0;
  assign pp_0_1_0 = pp_0_1;
  assign pp_0_1_1 = pp_1_1;
  assign pp_0_2_0 = pp_0_2;
  assign pp_0_2_1 = pp_1_2;
  assign pp_0_2_2 = pp_2_2;
  assign pp_0_3_0 = pp_0_3;
  assign pp_0_3_1 = pp_1_3;
  assign pp_0_3_2 = pp_2_3;
  assign pp_0_3_3 = pp_3_3;
  assign pp_0_4_0 = pp_0_4;
  assign pp_0_4_1 = pp_1_4;
  assign pp_0_4_2 = pp_2_4;
  assign pp_0_4_3 = pp_3_4;
  assign pp_0_4_4 = pp_4_4;
  assign pp_0_5_0 = pp_0_5;
  assign pp_0_5_1 = pp_1_5;
  assign pp_0_5_2 = pp_2_5;
  assign pp_0_5_3 = pp_3_5;
  assign pp_0_5_4 = pp_4_5;
  assign pp_0_5_5 = pp_5_5;
  assign pp_0_6_0 = pp_0_6;
  assign pp_0_6_1 = pp_1_6;
  assign pp_0_6_2 = pp_2_6;
  assign pp_0_6_3 = pp_3_6;
  assign pp_0_6_4 = pp_4_6;
  assign pp_0_6_5 = pp_5_6;
  assign pp_0_6_6 = pp_6_6;
  assign pp_0_7_0 = pp_0_7;
  assign pp_0_7_1 = pp_1_7;
  assign pp_0_7_2 = pp_2_7;
  assign pp_0_7_3 = pp_3_7;
  assign pp_0_7_4 = pp_4_7;
  assign pp_0_7_5 = pp_5_7;
  assign pp_0_7_6 = pp_6_7;
  assign pp_0_7_7 = pp_7_7;
  assign pp_0_8_0 = pp_0_8;
  assign pp_0_8_1 = pp_1_8;
  assign pp_0_8_2 = pp_2_8;
  assign pp_0_8_3 = pp_3_8;
  assign pp_0_8_4 = pp_4_8;
  assign pp_0_8_5 = pp_5_8;
  assign pp_0_8_6 = pp_6_8;
  assign pp_0_8_7 = pp_7_8;
  assign pp_0_8_8 = pp_8_8;
  assign pp_0_9_0 = pp_0_9;
  assign pp_0_9_1 = pp_1_9;
  assign pp_0_9_2 = pp_2_9;
  assign pp_0_9_3 = pp_3_9;
  assign pp_0_9_4 = pp_4_9;
  assign pp_0_9_5 = pp_5_9;
  assign pp_0_9_6 = pp_6_9;
  assign pp_0_9_7 = pp_7_9;
  assign pp_0_9_8 = pp_8_9;
  assign pp_0_9_9 = pp_9_9;
  assign pp_0_10_0 = pp_0_10;
  assign pp_0_10_1 = pp_1_10;
  assign pp_0_10_2 = pp_2_10;
  assign pp_0_10_3 = pp_3_10;
  assign pp_0_10_4 = pp_4_10;
  assign pp_0_10_5 = pp_5_10;
  assign pp_0_10_6 = pp_6_10;
  assign pp_0_10_7 = pp_7_10;
  assign pp_0_10_8 = pp_8_10;
  assign pp_0_10_9 = pp_9_10;
  assign pp_0_10_10 = pp_10_10;
  assign pp_0_11_0 = pp_0_11;
  assign pp_0_11_1 = pp_1_11;
  assign pp_0_11_2 = pp_2_11;
  assign pp_0_11_3 = pp_3_11;
  assign pp_0_11_4 = pp_4_11;
  assign pp_0_11_5 = pp_5_11;
  assign pp_0_11_6 = pp_6_11;
  assign pp_0_11_7 = pp_7_11;
  assign pp_0_11_8 = pp_8_11;
  assign pp_0_11_9 = pp_9_11;
  assign pp_0_11_10 = pp_10_11;
  assign pp_0_11_11 = pp_11_11;
  assign pp_0_12_0 = pp_0_12;
  assign pp_0_12_1 = pp_1_12;
  assign pp_0_12_2 = pp_2_12;
  assign pp_0_12_3 = pp_3_12;
  assign pp_0_12_4 = pp_4_12;
  assign pp_0_12_5 = pp_5_12;
  assign pp_0_12_6 = pp_6_12;
  assign pp_0_12_7 = pp_7_12;
  assign pp_0_12_8 = pp_8_12;
  assign pp_0_12_9 = pp_9_12;
  assign pp_0_12_10 = pp_10_12;
  assign pp_0_12_11 = pp_11_12;
  assign pp_0_12_12 = pp_12_12;
  assign pp_0_13_0 = pp_0_13;
  assign pp_0_13_1 = pp_1_13;
  assign pp_0_13_2 = pp_2_13;
  assign pp_0_13_3 = pp_3_13;
  assign pp_0_13_4 = pp_4_13;
  assign pp_0_13_5 = pp_5_13;
  assign pp_0_13_6 = pp_6_13;
  assign pp_0_13_7 = pp_7_13;
  assign pp_0_13_8 = pp_8_13;
  assign pp_0_13_9 = pp_9_13;
  assign pp_0_13_10 = pp_10_13;
  assign pp_0_13_11 = pp_11_13;
  assign pp_0_13_12 = pp_12_13;
  assign pp_0_13_13 = pp_13_13;
  assign pp_0_14_0 = pp_0_14;
  assign pp_0_14_1 = pp_1_14;
  assign pp_0_14_2 = pp_2_14;
  assign pp_0_14_3 = pp_3_14;
  assign pp_0_14_4 = pp_4_14;
  assign pp_0_14_5 = pp_5_14;
  assign pp_0_14_6 = pp_6_14;
  assign pp_0_14_7 = pp_7_14;
  assign pp_0_14_8 = pp_8_14;
  assign pp_0_14_9 = pp_9_14;
  assign pp_0_14_10 = pp_10_14;
  assign pp_0_14_11 = pp_11_14;
  assign pp_0_14_12 = pp_12_14;
  assign pp_0_14_13 = pp_13_14;
  assign pp_0_14_14 = pp_14_14;
  assign pp_0_15_0 = pp_0_15;
  assign pp_0_15_1 = pp_1_15;
  assign pp_0_15_2 = pp_2_15;
  assign pp_0_15_3 = pp_3_15;
  assign pp_0_15_4 = pp_4_15;
  assign pp_0_15_5 = pp_5_15;
  assign pp_0_15_6 = pp_6_15;
  assign pp_0_15_7 = pp_7_15;
  assign pp_0_15_8 = pp_8_15;
  assign pp_0_15_9 = pp_9_15;
  assign pp_0_15_10 = pp_10_15;
  assign pp_0_15_11 = pp_11_15;
  assign pp_0_15_12 = pp_12_15;
  assign pp_0_15_13 = pp_13_15;
  assign pp_0_15_14 = pp_14_15;
  assign pp_0_15_15 = pp_15_15;
  assign pp_0_16_0 = pp_0_16;
  assign pp_0_16_1 = pp_1_16;
  assign pp_0_16_2 = pp_2_16;
  assign pp_0_16_3 = pp_3_16;
  assign pp_0_16_4 = pp_4_16;
  assign pp_0_16_5 = pp_5_16;
  assign pp_0_16_6 = pp_6_16;
  assign pp_0_16_7 = pp_7_16;
  assign pp_0_16_8 = pp_8_16;
  assign pp_0_16_9 = pp_9_16;
  assign pp_0_16_10 = pp_10_16;
  assign pp_0_16_11 = pp_11_16;
  assign pp_0_16_12 = pp_12_16;
  assign pp_0_16_13 = pp_13_16;
  assign pp_0_16_14 = pp_14_16;
  assign pp_0_16_15 = pp_15_16;
  assign pp_0_16_16 = pp_16_16;
  assign pp_0_17_0 = pp_0_17;
  assign pp_0_17_1 = pp_1_17;
  assign pp_0_17_2 = pp_2_17;
  assign pp_0_17_3 = pp_3_17;
  assign pp_0_17_4 = pp_4_17;
  assign pp_0_17_5 = pp_5_17;
  assign pp_0_17_6 = pp_6_17;
  assign pp_0_17_7 = pp_7_17;
  assign pp_0_17_8 = pp_8_17;
  assign pp_0_17_9 = pp_9_17;
  assign pp_0_17_10 = pp_10_17;
  assign pp_0_17_11 = pp_11_17;
  assign pp_0_17_12 = pp_12_17;
  assign pp_0_17_13 = pp_13_17;
  assign pp_0_17_14 = pp_14_17;
  assign pp_0_17_15 = pp_15_17;
  assign pp_0_17_16 = pp_16_17;
  assign pp_0_17_17 = pp_17_17;
  assign pp_0_18_0 = pp_0_18;
  assign pp_0_18_1 = pp_1_18;
  assign pp_0_18_2 = pp_2_18;
  assign pp_0_18_3 = pp_3_18;
  assign pp_0_18_4 = pp_4_18;
  assign pp_0_18_5 = pp_5_18;
  assign pp_0_18_6 = pp_6_18;
  assign pp_0_18_7 = pp_7_18;
  assign pp_0_18_8 = pp_8_18;
  assign pp_0_18_9 = pp_9_18;
  assign pp_0_18_10 = pp_10_18;
  assign pp_0_18_11 = pp_11_18;
  assign pp_0_18_12 = pp_12_18;
  assign pp_0_18_13 = pp_13_18;
  assign pp_0_18_14 = pp_14_18;
  assign pp_0_18_15 = pp_15_18;
  assign pp_0_18_16 = pp_16_18;
  assign pp_0_18_17 = pp_17_18;
  assign pp_0_18_18 = pp_18_18;
  assign pp_0_19_0 = pp_0_19;
  assign pp_0_19_1 = pp_1_19;
  assign pp_0_19_2 = pp_2_19;
  assign pp_0_19_3 = pp_3_19;
  assign pp_0_19_4 = pp_4_19;
  assign pp_0_19_5 = pp_5_19;
  assign pp_0_19_6 = pp_6_19;
  assign pp_0_19_7 = pp_7_19;
  assign pp_0_19_8 = pp_8_19;
  assign pp_0_19_9 = pp_9_19;
  assign pp_0_19_10 = pp_10_19;
  assign pp_0_19_11 = pp_11_19;
  assign pp_0_19_12 = pp_12_19;
  assign pp_0_19_13 = pp_13_19;
  assign pp_0_19_14 = pp_14_19;
  assign pp_0_19_15 = pp_15_19;
  assign pp_0_19_16 = pp_16_19;
  assign pp_0_19_17 = pp_17_19;
  assign pp_0_19_18 = pp_18_19;
  assign pp_0_19_19 = pp_19_19;
  assign pp_0_20_0 = pp_0_20;
  assign pp_0_20_1 = pp_1_20;
  assign pp_0_20_2 = pp_2_20;
  assign pp_0_20_3 = pp_3_20;
  assign pp_0_20_4 = pp_4_20;
  assign pp_0_20_5 = pp_5_20;
  assign pp_0_20_6 = pp_6_20;
  assign pp_0_20_7 = pp_7_20;
  assign pp_0_20_8 = pp_8_20;
  assign pp_0_20_9 = pp_9_20;
  assign pp_0_20_10 = pp_10_20;
  assign pp_0_20_11 = pp_11_20;
  assign pp_0_20_12 = pp_12_20;
  assign pp_0_20_13 = pp_13_20;
  assign pp_0_20_14 = pp_14_20;
  assign pp_0_20_15 = pp_15_20;
  assign pp_0_20_16 = pp_16_20;
  assign pp_0_20_17 = pp_17_20;
  assign pp_0_20_18 = pp_18_20;
  assign pp_0_20_19 = pp_19_20;
  assign pp_0_20_20 = pp_20_20;
  assign pp_0_21_0 = pp_0_21;
  assign pp_0_21_1 = pp_1_21;
  assign pp_0_21_2 = pp_2_21;
  assign pp_0_21_3 = pp_3_21;
  assign pp_0_21_4 = pp_4_21;
  assign pp_0_21_5 = pp_5_21;
  assign pp_0_21_6 = pp_6_21;
  assign pp_0_21_7 = pp_7_21;
  assign pp_0_21_8 = pp_8_21;
  assign pp_0_21_9 = pp_9_21;
  assign pp_0_21_10 = pp_10_21;
  assign pp_0_21_11 = pp_11_21;
  assign pp_0_21_12 = pp_12_21;
  assign pp_0_21_13 = pp_13_21;
  assign pp_0_21_14 = pp_14_21;
  assign pp_0_21_15 = pp_15_21;
  assign pp_0_21_16 = pp_16_21;
  assign pp_0_21_17 = pp_17_21;
  assign pp_0_21_18 = pp_18_21;
  assign pp_0_21_19 = pp_19_21;
  assign pp_0_21_20 = pp_20_21;
  assign pp_0_21_21 = pp_21_21;
  assign pp_0_22_0 = pp_0_22;
  assign pp_0_22_1 = pp_1_22;
  assign pp_0_22_2 = pp_2_22;
  assign pp_0_22_3 = pp_3_22;
  assign pp_0_22_4 = pp_4_22;
  assign pp_0_22_5 = pp_5_22;
  assign pp_0_22_6 = pp_6_22;
  assign pp_0_22_7 = pp_7_22;
  assign pp_0_22_8 = pp_8_22;
  assign pp_0_22_9 = pp_9_22;
  assign pp_0_22_10 = pp_10_22;
  assign pp_0_22_11 = pp_11_22;
  assign pp_0_22_12 = pp_12_22;
  assign pp_0_22_13 = pp_13_22;
  assign pp_0_22_14 = pp_14_22;
  assign pp_0_22_15 = pp_15_22;
  assign pp_0_22_16 = pp_16_22;
  assign pp_0_22_17 = pp_17_22;
  assign pp_0_22_18 = pp_18_22;
  assign pp_0_22_19 = pp_19_22;
  assign pp_0_22_20 = pp_20_22;
  assign pp_0_22_21 = pp_21_22;
  assign pp_0_22_22 = pp_22_22;
  assign pp_0_23_0 = pp_0_23;
  assign pp_0_23_1 = pp_1_23;
  assign pp_0_23_2 = pp_2_23;
  assign pp_0_23_3 = pp_3_23;
  assign pp_0_23_4 = pp_4_23;
  assign pp_0_23_5 = pp_5_23;
  assign pp_0_23_6 = pp_6_23;
  assign pp_0_23_7 = pp_7_23;
  assign pp_0_23_8 = pp_8_23;
  assign pp_0_23_9 = pp_9_23;
  assign pp_0_23_10 = pp_10_23;
  assign pp_0_23_11 = pp_11_23;
  assign pp_0_23_12 = pp_12_23;
  assign pp_0_23_13 = pp_13_23;
  assign pp_0_23_14 = pp_14_23;
  assign pp_0_23_15 = pp_15_23;
  assign pp_0_23_16 = pp_16_23;
  assign pp_0_23_17 = pp_17_23;
  assign pp_0_23_18 = pp_18_23;
  assign pp_0_23_19 = pp_19_23;
  assign pp_0_23_20 = pp_20_23;
  assign pp_0_23_21 = pp_21_23;
  assign pp_0_23_22 = pp_22_23;
  assign pp_0_23_23 = pp_23_23;
  assign pp_0_24_0 = pp_0_24;
  assign pp_0_24_1 = pp_1_24;
  assign pp_0_24_2 = pp_2_24;
  assign pp_0_24_3 = pp_3_24;
  assign pp_0_24_4 = pp_4_24;
  assign pp_0_24_5 = pp_5_24;
  assign pp_0_24_6 = pp_6_24;
  assign pp_0_24_7 = pp_7_24;
  assign pp_0_24_8 = pp_8_24;
  assign pp_0_24_9 = pp_9_24;
  assign pp_0_24_10 = pp_10_24;
  assign pp_0_24_11 = pp_11_24;
  assign pp_0_24_12 = pp_12_24;
  assign pp_0_24_13 = pp_13_24;
  assign pp_0_24_14 = pp_14_24;
  assign pp_0_24_15 = pp_15_24;
  assign pp_0_24_16 = pp_16_24;
  assign pp_0_24_17 = pp_17_24;
  assign pp_0_24_18 = pp_18_24;
  assign pp_0_24_19 = pp_19_24;
  assign pp_0_24_20 = pp_20_24;
  assign pp_0_24_21 = pp_21_24;
  assign pp_0_24_22 = pp_22_24;
  assign pp_0_24_23 = pp_23_24;
  assign pp_0_24_24 = pp_24_24;
  assign pp_0_25_0 = pp_0_25;
  assign pp_0_25_1 = pp_1_25;
  assign pp_0_25_2 = pp_2_25;
  assign pp_0_25_3 = pp_3_25;
  assign pp_0_25_4 = pp_4_25;
  assign pp_0_25_5 = pp_5_25;
  assign pp_0_25_6 = pp_6_25;
  assign pp_0_25_7 = pp_7_25;
  assign pp_0_25_8 = pp_8_25;
  assign pp_0_25_9 = pp_9_25;
  assign pp_0_25_10 = pp_10_25;
  assign pp_0_25_11 = pp_11_25;
  assign pp_0_25_12 = pp_12_25;
  assign pp_0_25_13 = pp_13_25;
  assign pp_0_25_14 = pp_14_25;
  assign pp_0_25_15 = pp_15_25;
  assign pp_0_25_16 = pp_16_25;
  assign pp_0_25_17 = pp_17_25;
  assign pp_0_25_18 = pp_18_25;
  assign pp_0_25_19 = pp_19_25;
  assign pp_0_25_20 = pp_20_25;
  assign pp_0_25_21 = pp_21_25;
  assign pp_0_25_22 = pp_22_25;
  assign pp_0_25_23 = pp_23_25;
  assign pp_0_25_24 = pp_24_25;
  assign pp_0_25_25 = pp_25_25;
  assign pp_0_26_0 = pp_0_26;
  assign pp_0_26_1 = pp_1_26;
  assign pp_0_26_2 = pp_2_26;
  assign pp_0_26_3 = pp_3_26;
  assign pp_0_26_4 = pp_4_26;
  assign pp_0_26_5 = pp_5_26;
  assign pp_0_26_6 = pp_6_26;
  assign pp_0_26_7 = pp_7_26;
  assign pp_0_26_8 = pp_8_26;
  assign pp_0_26_9 = pp_9_26;
  assign pp_0_26_10 = pp_10_26;
  assign pp_0_26_11 = pp_11_26;
  assign pp_0_26_12 = pp_12_26;
  assign pp_0_26_13 = pp_13_26;
  assign pp_0_26_14 = pp_14_26;
  assign pp_0_26_15 = pp_15_26;
  assign pp_0_26_16 = pp_16_26;
  assign pp_0_26_17 = pp_17_26;
  assign pp_0_26_18 = pp_18_26;
  assign pp_0_26_19 = pp_19_26;
  assign pp_0_26_20 = pp_20_26;
  assign pp_0_26_21 = pp_21_26;
  assign pp_0_26_22 = pp_22_26;
  assign pp_0_26_23 = pp_23_26;
  assign pp_0_26_24 = pp_24_26;
  assign pp_0_26_25 = pp_25_26;
  assign pp_0_26_26 = pp_26_26;
  assign pp_0_27_0 = pp_0_27;
  assign pp_0_27_1 = pp_1_27;
  assign pp_0_27_2 = pp_2_27;
  assign pp_0_27_3 = pp_3_27;
  assign pp_0_27_4 = pp_4_27;
  assign pp_0_27_5 = pp_5_27;
  assign pp_0_27_6 = pp_6_27;
  assign pp_0_27_7 = pp_7_27;
  assign pp_0_27_8 = pp_8_27;
  assign pp_0_27_9 = pp_9_27;
  assign pp_0_27_10 = pp_10_27;
  assign pp_0_27_11 = pp_11_27;
  assign pp_0_27_12 = pp_12_27;
  assign pp_0_27_13 = pp_13_27;
  assign pp_0_27_14 = pp_14_27;
  assign pp_0_27_15 = pp_15_27;
  assign pp_0_27_16 = pp_16_27;
  assign pp_0_27_17 = pp_17_27;
  assign pp_0_27_18 = pp_18_27;
  assign pp_0_27_19 = pp_19_27;
  assign pp_0_27_20 = pp_20_27;
  assign pp_0_27_21 = pp_21_27;
  assign pp_0_27_22 = pp_22_27;
  assign pp_0_27_23 = pp_23_27;
  assign pp_0_27_24 = pp_24_27;
  assign pp_0_27_25 = pp_25_27;
  assign pp_0_27_26 = pp_26_27;
  assign pp_0_27_27 = pp_27_27;
  assign pp_0_28_0 = pp_0_28;
  assign pp_0_28_1 = pp_1_28;
  assign pp_0_28_2 = pp_2_28;
  assign pp_0_28_3 = pp_3_28;
  assign pp_0_28_4 = pp_4_28;
  assign pp_0_28_5 = pp_5_28;
  assign pp_0_28_6 = pp_6_28;
  assign pp_0_28_7 = pp_7_28;
  assign pp_0_28_8 = pp_8_28;
  assign pp_0_28_9 = pp_9_28;
  assign pp_0_28_10 = pp_10_28;
  assign pp_0_28_11 = pp_11_28;
  assign pp_0_28_12 = pp_12_28;
  assign pp_0_28_13 = pp_13_28;
  assign pp_0_28_14 = pp_14_28;
  assign pp_0_28_15 = pp_15_28;
  assign pp_0_28_16 = pp_16_28;
  assign pp_0_28_17 = pp_17_28;
  assign pp_0_28_18 = pp_18_28;
  assign pp_0_28_19 = pp_19_28;
  assign pp_0_28_20 = pp_20_28;
  assign pp_0_28_21 = pp_21_28;
  assign pp_0_28_22 = pp_22_28;
  assign pp_0_28_23 = pp_23_28;
  assign pp_0_28_24 = pp_24_28;
  assign pp_0_28_25 = pp_25_28;
  assign pp_0_28_26 = pp_26_28;
  assign pp_0_28_27 = pp_27_28;
  assign pp_0_28_28 = pp_28_28;
  assign pp_0_29_0 = pp_0_29;
  assign pp_0_29_1 = pp_1_29;
  assign pp_0_29_2 = pp_2_29;
  assign pp_0_29_3 = pp_3_29;
  assign pp_0_29_4 = pp_4_29;
  assign pp_0_29_5 = pp_5_29;
  assign pp_0_29_6 = pp_6_29;
  assign pp_0_29_7 = pp_7_29;
  assign pp_0_29_8 = pp_8_29;
  assign pp_0_29_9 = pp_9_29;
  assign pp_0_29_10 = pp_10_29;
  assign pp_0_29_11 = pp_11_29;
  assign pp_0_29_12 = pp_12_29;
  assign pp_0_29_13 = pp_13_29;
  assign pp_0_29_14 = pp_14_29;
  assign pp_0_29_15 = pp_15_29;
  assign pp_0_29_16 = pp_16_29;
  assign pp_0_29_17 = pp_17_29;
  assign pp_0_29_18 = pp_18_29;
  assign pp_0_29_19 = pp_19_29;
  assign pp_0_29_20 = pp_20_29;
  assign pp_0_29_21 = pp_21_29;
  assign pp_0_29_22 = pp_22_29;
  assign pp_0_29_23 = pp_23_29;
  assign pp_0_29_24 = pp_24_29;
  assign pp_0_29_25 = pp_25_29;
  assign pp_0_29_26 = pp_26_29;
  assign pp_0_29_27 = pp_27_29;
  assign pp_0_29_28 = pp_28_29;
  assign pp_0_29_29 = pp_29_29;
  assign pp_0_30_0 = pp_0_30;
  assign pp_0_30_1 = pp_1_30;
  assign pp_0_30_2 = pp_2_30;
  assign pp_0_30_3 = pp_3_30;
  assign pp_0_30_4 = pp_4_30;
  assign pp_0_30_5 = pp_5_30;
  assign pp_0_30_6 = pp_6_30;
  assign pp_0_30_7 = pp_7_30;
  assign pp_0_30_8 = pp_8_30;
  assign pp_0_30_9 = pp_9_30;
  assign pp_0_30_10 = pp_10_30;
  assign pp_0_30_11 = pp_11_30;
  assign pp_0_30_12 = pp_12_30;
  assign pp_0_30_13 = pp_13_30;
  assign pp_0_30_14 = pp_14_30;
  assign pp_0_30_15 = pp_15_30;
  assign pp_0_30_16 = pp_16_30;
  assign pp_0_30_17 = pp_17_30;
  assign pp_0_30_18 = pp_18_30;
  assign pp_0_30_19 = pp_19_30;
  assign pp_0_30_20 = pp_20_30;
  assign pp_0_30_21 = pp_21_30;
  assign pp_0_30_22 = pp_22_30;
  assign pp_0_30_23 = pp_23_30;
  assign pp_0_30_24 = pp_24_30;
  assign pp_0_30_25 = pp_25_30;
  assign pp_0_30_26 = pp_26_30;
  assign pp_0_30_27 = pp_27_30;
  assign pp_0_30_28 = pp_28_30;
  assign pp_0_30_29 = pp_29_30;
  assign pp_0_30_30 = pp_30_30;
  assign pp_0_31_0 = pp_0_31;
  assign pp_0_31_1 = pp_1_31;
  assign pp_0_31_2 = pp_2_31;
  assign pp_0_31_3 = pp_3_31;
  assign pp_0_31_4 = pp_4_31;
  assign pp_0_31_5 = pp_5_31;
  assign pp_0_31_6 = pp_6_31;
  assign pp_0_31_7 = pp_7_31;
  assign pp_0_31_8 = pp_8_31;
  assign pp_0_31_9 = pp_9_31;
  assign pp_0_31_10 = pp_10_31;
  assign pp_0_31_11 = pp_11_31;
  assign pp_0_31_12 = pp_12_31;
  assign pp_0_31_13 = pp_13_31;
  assign pp_0_31_14 = pp_14_31;
  assign pp_0_31_15 = pp_15_31;
  assign pp_0_31_16 = pp_16_31;
  assign pp_0_31_17 = pp_17_31;
  assign pp_0_31_18 = pp_18_31;
  assign pp_0_31_19 = pp_19_31;
  assign pp_0_31_20 = pp_20_31;
  assign pp_0_31_21 = pp_21_31;
  assign pp_0_31_22 = pp_22_31;
  assign pp_0_31_23 = pp_23_31;
  assign pp_0_31_24 = pp_24_31;
  assign pp_0_31_25 = pp_25_31;
  assign pp_0_31_26 = pp_26_31;
  assign pp_0_31_27 = pp_27_31;
  assign pp_0_31_28 = pp_28_31;
  assign pp_0_31_29 = pp_29_31;
  assign pp_0_31_30 = pp_30_31;
  assign pp_0_31_31 = pp_31_31;
  assign pp_0_32_0 = pp_1_32;
  assign pp_0_32_1 = pp_2_32;
  assign pp_0_32_2 = pp_3_32;
  assign pp_0_32_3 = pp_4_32;
  assign pp_0_32_4 = pp_5_32;
  assign pp_0_32_5 = pp_6_32;
  assign pp_0_32_6 = pp_7_32;
  assign pp_0_32_7 = pp_8_32;
  assign pp_0_32_8 = pp_9_32;
  assign pp_0_32_9 = pp_10_32;
  assign pp_0_32_10 = pp_11_32;
  assign pp_0_32_11 = pp_12_32;
  assign pp_0_32_12 = pp_13_32;
  assign pp_0_32_13 = pp_14_32;
  assign pp_0_32_14 = pp_15_32;
  assign pp_0_32_15 = pp_16_32;
  assign pp_0_32_16 = pp_17_32;
  assign pp_0_32_17 = pp_18_32;
  assign pp_0_32_18 = pp_19_32;
  assign pp_0_32_19 = pp_20_32;
  assign pp_0_32_20 = pp_21_32;
  assign pp_0_32_21 = pp_22_32;
  assign pp_0_32_22 = pp_23_32;
  assign pp_0_32_23 = pp_24_32;
  assign pp_0_32_24 = pp_25_32;
  assign pp_0_32_25 = pp_26_32;
  assign pp_0_32_26 = pp_27_32;
  assign pp_0_32_27 = pp_28_32;
  assign pp_0_32_28 = pp_29_32;
  assign pp_0_32_29 = pp_30_32;
  assign pp_0_32_30 = pp_31_32;
  assign pp_0_33_0 = pp_2_33;
  assign pp_0_33_1 = pp_3_33;
  assign pp_0_33_2 = pp_4_33;
  assign pp_0_33_3 = pp_5_33;
  assign pp_0_33_4 = pp_6_33;
  assign pp_0_33_5 = pp_7_33;
  assign pp_0_33_6 = pp_8_33;
  assign pp_0_33_7 = pp_9_33;
  assign pp_0_33_8 = pp_10_33;
  assign pp_0_33_9 = pp_11_33;
  assign pp_0_33_10 = pp_12_33;
  assign pp_0_33_11 = pp_13_33;
  assign pp_0_33_12 = pp_14_33;
  assign pp_0_33_13 = pp_15_33;
  assign pp_0_33_14 = pp_16_33;
  assign pp_0_33_15 = pp_17_33;
  assign pp_0_33_16 = pp_18_33;
  assign pp_0_33_17 = pp_19_33;
  assign pp_0_33_18 = pp_20_33;
  assign pp_0_33_19 = pp_21_33;
  assign pp_0_33_20 = pp_22_33;
  assign pp_0_33_21 = pp_23_33;
  assign pp_0_33_22 = pp_24_33;
  assign pp_0_33_23 = pp_25_33;
  assign pp_0_33_24 = pp_26_33;
  assign pp_0_33_25 = pp_27_33;
  assign pp_0_33_26 = pp_28_33;
  assign pp_0_33_27 = pp_29_33;
  assign pp_0_33_28 = pp_30_33;
  assign pp_0_33_29 = pp_31_33;
  assign pp_0_34_0 = pp_3_34;
  assign pp_0_34_1 = pp_4_34;
  assign pp_0_34_2 = pp_5_34;
  assign pp_0_34_3 = pp_6_34;
  assign pp_0_34_4 = pp_7_34;
  assign pp_0_34_5 = pp_8_34;
  assign pp_0_34_6 = pp_9_34;
  assign pp_0_34_7 = pp_10_34;
  assign pp_0_34_8 = pp_11_34;
  assign pp_0_34_9 = pp_12_34;
  assign pp_0_34_10 = pp_13_34;
  assign pp_0_34_11 = pp_14_34;
  assign pp_0_34_12 = pp_15_34;
  assign pp_0_34_13 = pp_16_34;
  assign pp_0_34_14 = pp_17_34;
  assign pp_0_34_15 = pp_18_34;
  assign pp_0_34_16 = pp_19_34;
  assign pp_0_34_17 = pp_20_34;
  assign pp_0_34_18 = pp_21_34;
  assign pp_0_34_19 = pp_22_34;
  assign pp_0_34_20 = pp_23_34;
  assign pp_0_34_21 = pp_24_34;
  assign pp_0_34_22 = pp_25_34;
  assign pp_0_34_23 = pp_26_34;
  assign pp_0_34_24 = pp_27_34;
  assign pp_0_34_25 = pp_28_34;
  assign pp_0_34_26 = pp_29_34;
  assign pp_0_34_27 = pp_30_34;
  assign pp_0_34_28 = pp_31_34;
  assign pp_0_35_0 = pp_4_35;
  assign pp_0_35_1 = pp_5_35;
  assign pp_0_35_2 = pp_6_35;
  assign pp_0_35_3 = pp_7_35;
  assign pp_0_35_4 = pp_8_35;
  assign pp_0_35_5 = pp_9_35;
  assign pp_0_35_6 = pp_10_35;
  assign pp_0_35_7 = pp_11_35;
  assign pp_0_35_8 = pp_12_35;
  assign pp_0_35_9 = pp_13_35;
  assign pp_0_35_10 = pp_14_35;
  assign pp_0_35_11 = pp_15_35;
  assign pp_0_35_12 = pp_16_35;
  assign pp_0_35_13 = pp_17_35;
  assign pp_0_35_14 = pp_18_35;
  assign pp_0_35_15 = pp_19_35;
  assign pp_0_35_16 = pp_20_35;
  assign pp_0_35_17 = pp_21_35;
  assign pp_0_35_18 = pp_22_35;
  assign pp_0_35_19 = pp_23_35;
  assign pp_0_35_20 = pp_24_35;
  assign pp_0_35_21 = pp_25_35;
  assign pp_0_35_22 = pp_26_35;
  assign pp_0_35_23 = pp_27_35;
  assign pp_0_35_24 = pp_28_35;
  assign pp_0_35_25 = pp_29_35;
  assign pp_0_35_26 = pp_30_35;
  assign pp_0_35_27 = pp_31_35;
  assign pp_0_36_0 = pp_5_36;
  assign pp_0_36_1 = pp_6_36;
  assign pp_0_36_2 = pp_7_36;
  assign pp_0_36_3 = pp_8_36;
  assign pp_0_36_4 = pp_9_36;
  assign pp_0_36_5 = pp_10_36;
  assign pp_0_36_6 = pp_11_36;
  assign pp_0_36_7 = pp_12_36;
  assign pp_0_36_8 = pp_13_36;
  assign pp_0_36_9 = pp_14_36;
  assign pp_0_36_10 = pp_15_36;
  assign pp_0_36_11 = pp_16_36;
  assign pp_0_36_12 = pp_17_36;
  assign pp_0_36_13 = pp_18_36;
  assign pp_0_36_14 = pp_19_36;
  assign pp_0_36_15 = pp_20_36;
  assign pp_0_36_16 = pp_21_36;
  assign pp_0_36_17 = pp_22_36;
  assign pp_0_36_18 = pp_23_36;
  assign pp_0_36_19 = pp_24_36;
  assign pp_0_36_20 = pp_25_36;
  assign pp_0_36_21 = pp_26_36;
  assign pp_0_36_22 = pp_27_36;
  assign pp_0_36_23 = pp_28_36;
  assign pp_0_36_24 = pp_29_36;
  assign pp_0_36_25 = pp_30_36;
  assign pp_0_36_26 = pp_31_36;
  assign pp_0_37_0 = pp_6_37;
  assign pp_0_37_1 = pp_7_37;
  assign pp_0_37_2 = pp_8_37;
  assign pp_0_37_3 = pp_9_37;
  assign pp_0_37_4 = pp_10_37;
  assign pp_0_37_5 = pp_11_37;
  assign pp_0_37_6 = pp_12_37;
  assign pp_0_37_7 = pp_13_37;
  assign pp_0_37_8 = pp_14_37;
  assign pp_0_37_9 = pp_15_37;
  assign pp_0_37_10 = pp_16_37;
  assign pp_0_37_11 = pp_17_37;
  assign pp_0_37_12 = pp_18_37;
  assign pp_0_37_13 = pp_19_37;
  assign pp_0_37_14 = pp_20_37;
  assign pp_0_37_15 = pp_21_37;
  assign pp_0_37_16 = pp_22_37;
  assign pp_0_37_17 = pp_23_37;
  assign pp_0_37_18 = pp_24_37;
  assign pp_0_37_19 = pp_25_37;
  assign pp_0_37_20 = pp_26_37;
  assign pp_0_37_21 = pp_27_37;
  assign pp_0_37_22 = pp_28_37;
  assign pp_0_37_23 = pp_29_37;
  assign pp_0_37_24 = pp_30_37;
  assign pp_0_37_25 = pp_31_37;
  assign pp_0_38_0 = pp_7_38;
  assign pp_0_38_1 = pp_8_38;
  assign pp_0_38_2 = pp_9_38;
  assign pp_0_38_3 = pp_10_38;
  assign pp_0_38_4 = pp_11_38;
  assign pp_0_38_5 = pp_12_38;
  assign pp_0_38_6 = pp_13_38;
  assign pp_0_38_7 = pp_14_38;
  assign pp_0_38_8 = pp_15_38;
  assign pp_0_38_9 = pp_16_38;
  assign pp_0_38_10 = pp_17_38;
  assign pp_0_38_11 = pp_18_38;
  assign pp_0_38_12 = pp_19_38;
  assign pp_0_38_13 = pp_20_38;
  assign pp_0_38_14 = pp_21_38;
  assign pp_0_38_15 = pp_22_38;
  assign pp_0_38_16 = pp_23_38;
  assign pp_0_38_17 = pp_24_38;
  assign pp_0_38_18 = pp_25_38;
  assign pp_0_38_19 = pp_26_38;
  assign pp_0_38_20 = pp_27_38;
  assign pp_0_38_21 = pp_28_38;
  assign pp_0_38_22 = pp_29_38;
  assign pp_0_38_23 = pp_30_38;
  assign pp_0_38_24 = pp_31_38;
  assign pp_0_39_0 = pp_8_39;
  assign pp_0_39_1 = pp_9_39;
  assign pp_0_39_2 = pp_10_39;
  assign pp_0_39_3 = pp_11_39;
  assign pp_0_39_4 = pp_12_39;
  assign pp_0_39_5 = pp_13_39;
  assign pp_0_39_6 = pp_14_39;
  assign pp_0_39_7 = pp_15_39;
  assign pp_0_39_8 = pp_16_39;
  assign pp_0_39_9 = pp_17_39;
  assign pp_0_39_10 = pp_18_39;
  assign pp_0_39_11 = pp_19_39;
  assign pp_0_39_12 = pp_20_39;
  assign pp_0_39_13 = pp_21_39;
  assign pp_0_39_14 = pp_22_39;
  assign pp_0_39_15 = pp_23_39;
  assign pp_0_39_16 = pp_24_39;
  assign pp_0_39_17 = pp_25_39;
  assign pp_0_39_18 = pp_26_39;
  assign pp_0_39_19 = pp_27_39;
  assign pp_0_39_20 = pp_28_39;
  assign pp_0_39_21 = pp_29_39;
  assign pp_0_39_22 = pp_30_39;
  assign pp_0_39_23 = pp_31_39;
  assign pp_0_40_0 = pp_9_40;
  assign pp_0_40_1 = pp_10_40;
  assign pp_0_40_2 = pp_11_40;
  assign pp_0_40_3 = pp_12_40;
  assign pp_0_40_4 = pp_13_40;
  assign pp_0_40_5 = pp_14_40;
  assign pp_0_40_6 = pp_15_40;
  assign pp_0_40_7 = pp_16_40;
  assign pp_0_40_8 = pp_17_40;
  assign pp_0_40_9 = pp_18_40;
  assign pp_0_40_10 = pp_19_40;
  assign pp_0_40_11 = pp_20_40;
  assign pp_0_40_12 = pp_21_40;
  assign pp_0_40_13 = pp_22_40;
  assign pp_0_40_14 = pp_23_40;
  assign pp_0_40_15 = pp_24_40;
  assign pp_0_40_16 = pp_25_40;
  assign pp_0_40_17 = pp_26_40;
  assign pp_0_40_18 = pp_27_40;
  assign pp_0_40_19 = pp_28_40;
  assign pp_0_40_20 = pp_29_40;
  assign pp_0_40_21 = pp_30_40;
  assign pp_0_40_22 = pp_31_40;
  assign pp_0_41_0 = pp_10_41;
  assign pp_0_41_1 = pp_11_41;
  assign pp_0_41_2 = pp_12_41;
  assign pp_0_41_3 = pp_13_41;
  assign pp_0_41_4 = pp_14_41;
  assign pp_0_41_5 = pp_15_41;
  assign pp_0_41_6 = pp_16_41;
  assign pp_0_41_7 = pp_17_41;
  assign pp_0_41_8 = pp_18_41;
  assign pp_0_41_9 = pp_19_41;
  assign pp_0_41_10 = pp_20_41;
  assign pp_0_41_11 = pp_21_41;
  assign pp_0_41_12 = pp_22_41;
  assign pp_0_41_13 = pp_23_41;
  assign pp_0_41_14 = pp_24_41;
  assign pp_0_41_15 = pp_25_41;
  assign pp_0_41_16 = pp_26_41;
  assign pp_0_41_17 = pp_27_41;
  assign pp_0_41_18 = pp_28_41;
  assign pp_0_41_19 = pp_29_41;
  assign pp_0_41_20 = pp_30_41;
  assign pp_0_41_21 = pp_31_41;
  assign pp_0_42_0 = pp_11_42;
  assign pp_0_42_1 = pp_12_42;
  assign pp_0_42_2 = pp_13_42;
  assign pp_0_42_3 = pp_14_42;
  assign pp_0_42_4 = pp_15_42;
  assign pp_0_42_5 = pp_16_42;
  assign pp_0_42_6 = pp_17_42;
  assign pp_0_42_7 = pp_18_42;
  assign pp_0_42_8 = pp_19_42;
  assign pp_0_42_9 = pp_20_42;
  assign pp_0_42_10 = pp_21_42;
  assign pp_0_42_11 = pp_22_42;
  assign pp_0_42_12 = pp_23_42;
  assign pp_0_42_13 = pp_24_42;
  assign pp_0_42_14 = pp_25_42;
  assign pp_0_42_15 = pp_26_42;
  assign pp_0_42_16 = pp_27_42;
  assign pp_0_42_17 = pp_28_42;
  assign pp_0_42_18 = pp_29_42;
  assign pp_0_42_19 = pp_30_42;
  assign pp_0_42_20 = pp_31_42;
  assign pp_0_43_0 = pp_12_43;
  assign pp_0_43_1 = pp_13_43;
  assign pp_0_43_2 = pp_14_43;
  assign pp_0_43_3 = pp_15_43;
  assign pp_0_43_4 = pp_16_43;
  assign pp_0_43_5 = pp_17_43;
  assign pp_0_43_6 = pp_18_43;
  assign pp_0_43_7 = pp_19_43;
  assign pp_0_43_8 = pp_20_43;
  assign pp_0_43_9 = pp_21_43;
  assign pp_0_43_10 = pp_22_43;
  assign pp_0_43_11 = pp_23_43;
  assign pp_0_43_12 = pp_24_43;
  assign pp_0_43_13 = pp_25_43;
  assign pp_0_43_14 = pp_26_43;
  assign pp_0_43_15 = pp_27_43;
  assign pp_0_43_16 = pp_28_43;
  assign pp_0_43_17 = pp_29_43;
  assign pp_0_43_18 = pp_30_43;
  assign pp_0_43_19 = pp_31_43;
  assign pp_0_44_0 = pp_13_44;
  assign pp_0_44_1 = pp_14_44;
  assign pp_0_44_2 = pp_15_44;
  assign pp_0_44_3 = pp_16_44;
  assign pp_0_44_4 = pp_17_44;
  assign pp_0_44_5 = pp_18_44;
  assign pp_0_44_6 = pp_19_44;
  assign pp_0_44_7 = pp_20_44;
  assign pp_0_44_8 = pp_21_44;
  assign pp_0_44_9 = pp_22_44;
  assign pp_0_44_10 = pp_23_44;
  assign pp_0_44_11 = pp_24_44;
  assign pp_0_44_12 = pp_25_44;
  assign pp_0_44_13 = pp_26_44;
  assign pp_0_44_14 = pp_27_44;
  assign pp_0_44_15 = pp_28_44;
  assign pp_0_44_16 = pp_29_44;
  assign pp_0_44_17 = pp_30_44;
  assign pp_0_44_18 = pp_31_44;
  assign pp_0_45_0 = pp_14_45;
  assign pp_0_45_1 = pp_15_45;
  assign pp_0_45_2 = pp_16_45;
  assign pp_0_45_3 = pp_17_45;
  assign pp_0_45_4 = pp_18_45;
  assign pp_0_45_5 = pp_19_45;
  assign pp_0_45_6 = pp_20_45;
  assign pp_0_45_7 = pp_21_45;
  assign pp_0_45_8 = pp_22_45;
  assign pp_0_45_9 = pp_23_45;
  assign pp_0_45_10 = pp_24_45;
  assign pp_0_45_11 = pp_25_45;
  assign pp_0_45_12 = pp_26_45;
  assign pp_0_45_13 = pp_27_45;
  assign pp_0_45_14 = pp_28_45;
  assign pp_0_45_15 = pp_29_45;
  assign pp_0_45_16 = pp_30_45;
  assign pp_0_45_17 = pp_31_45;
  assign pp_0_46_0 = pp_15_46;
  assign pp_0_46_1 = pp_16_46;
  assign pp_0_46_2 = pp_17_46;
  assign pp_0_46_3 = pp_18_46;
  assign pp_0_46_4 = pp_19_46;
  assign pp_0_46_5 = pp_20_46;
  assign pp_0_46_6 = pp_21_46;
  assign pp_0_46_7 = pp_22_46;
  assign pp_0_46_8 = pp_23_46;
  assign pp_0_46_9 = pp_24_46;
  assign pp_0_46_10 = pp_25_46;
  assign pp_0_46_11 = pp_26_46;
  assign pp_0_46_12 = pp_27_46;
  assign pp_0_46_13 = pp_28_46;
  assign pp_0_46_14 = pp_29_46;
  assign pp_0_46_15 = pp_30_46;
  assign pp_0_46_16 = pp_31_46;
  assign pp_0_47_0 = pp_16_47;
  assign pp_0_47_1 = pp_17_47;
  assign pp_0_47_2 = pp_18_47;
  assign pp_0_47_3 = pp_19_47;
  assign pp_0_47_4 = pp_20_47;
  assign pp_0_47_5 = pp_21_47;
  assign pp_0_47_6 = pp_22_47;
  assign pp_0_47_7 = pp_23_47;
  assign pp_0_47_8 = pp_24_47;
  assign pp_0_47_9 = pp_25_47;
  assign pp_0_47_10 = pp_26_47;
  assign pp_0_47_11 = pp_27_47;
  assign pp_0_47_12 = pp_28_47;
  assign pp_0_47_13 = pp_29_47;
  assign pp_0_47_14 = pp_30_47;
  assign pp_0_47_15 = pp_31_47;
  assign pp_0_48_0 = pp_17_48;
  assign pp_0_48_1 = pp_18_48;
  assign pp_0_48_2 = pp_19_48;
  assign pp_0_48_3 = pp_20_48;
  assign pp_0_48_4 = pp_21_48;
  assign pp_0_48_5 = pp_22_48;
  assign pp_0_48_6 = pp_23_48;
  assign pp_0_48_7 = pp_24_48;
  assign pp_0_48_8 = pp_25_48;
  assign pp_0_48_9 = pp_26_48;
  assign pp_0_48_10 = pp_27_48;
  assign pp_0_48_11 = pp_28_48;
  assign pp_0_48_12 = pp_29_48;
  assign pp_0_48_13 = pp_30_48;
  assign pp_0_48_14 = pp_31_48;
  assign pp_0_49_0 = pp_18_49;
  assign pp_0_49_1 = pp_19_49;
  assign pp_0_49_2 = pp_20_49;
  assign pp_0_49_3 = pp_21_49;
  assign pp_0_49_4 = pp_22_49;
  assign pp_0_49_5 = pp_23_49;
  assign pp_0_49_6 = pp_24_49;
  assign pp_0_49_7 = pp_25_49;
  assign pp_0_49_8 = pp_26_49;
  assign pp_0_49_9 = pp_27_49;
  assign pp_0_49_10 = pp_28_49;
  assign pp_0_49_11 = pp_29_49;
  assign pp_0_49_12 = pp_30_49;
  assign pp_0_49_13 = pp_31_49;
  assign pp_0_50_0 = pp_19_50;
  assign pp_0_50_1 = pp_20_50;
  assign pp_0_50_2 = pp_21_50;
  assign pp_0_50_3 = pp_22_50;
  assign pp_0_50_4 = pp_23_50;
  assign pp_0_50_5 = pp_24_50;
  assign pp_0_50_6 = pp_25_50;
  assign pp_0_50_7 = pp_26_50;
  assign pp_0_50_8 = pp_27_50;
  assign pp_0_50_9 = pp_28_50;
  assign pp_0_50_10 = pp_29_50;
  assign pp_0_50_11 = pp_30_50;
  assign pp_0_50_12 = pp_31_50;
  assign pp_0_51_0 = pp_20_51;
  assign pp_0_51_1 = pp_21_51;
  assign pp_0_51_2 = pp_22_51;
  assign pp_0_51_3 = pp_23_51;
  assign pp_0_51_4 = pp_24_51;
  assign pp_0_51_5 = pp_25_51;
  assign pp_0_51_6 = pp_26_51;
  assign pp_0_51_7 = pp_27_51;
  assign pp_0_51_8 = pp_28_51;
  assign pp_0_51_9 = pp_29_51;
  assign pp_0_51_10 = pp_30_51;
  assign pp_0_51_11 = pp_31_51;
  assign pp_0_52_0 = pp_21_52;
  assign pp_0_52_1 = pp_22_52;
  assign pp_0_52_2 = pp_23_52;
  assign pp_0_52_3 = pp_24_52;
  assign pp_0_52_4 = pp_25_52;
  assign pp_0_52_5 = pp_26_52;
  assign pp_0_52_6 = pp_27_52;
  assign pp_0_52_7 = pp_28_52;
  assign pp_0_52_8 = pp_29_52;
  assign pp_0_52_9 = pp_30_52;
  assign pp_0_52_10 = pp_31_52;
  assign pp_0_53_0 = pp_22_53;
  assign pp_0_53_1 = pp_23_53;
  assign pp_0_53_2 = pp_24_53;
  assign pp_0_53_3 = pp_25_53;
  assign pp_0_53_4 = pp_26_53;
  assign pp_0_53_5 = pp_27_53;
  assign pp_0_53_6 = pp_28_53;
  assign pp_0_53_7 = pp_29_53;
  assign pp_0_53_8 = pp_30_53;
  assign pp_0_53_9 = pp_31_53;
  assign pp_0_54_0 = pp_23_54;
  assign pp_0_54_1 = pp_24_54;
  assign pp_0_54_2 = pp_25_54;
  assign pp_0_54_3 = pp_26_54;
  assign pp_0_54_4 = pp_27_54;
  assign pp_0_54_5 = pp_28_54;
  assign pp_0_54_6 = pp_29_54;
  assign pp_0_54_7 = pp_30_54;
  assign pp_0_54_8 = pp_31_54;
  assign pp_0_55_0 = pp_24_55;
  assign pp_0_55_1 = pp_25_55;
  assign pp_0_55_2 = pp_26_55;
  assign pp_0_55_3 = pp_27_55;
  assign pp_0_55_4 = pp_28_55;
  assign pp_0_55_5 = pp_29_55;
  assign pp_0_55_6 = pp_30_55;
  assign pp_0_55_7 = pp_31_55;
  assign pp_0_56_0 = pp_25_56;
  assign pp_0_56_1 = pp_26_56;
  assign pp_0_56_2 = pp_27_56;
  assign pp_0_56_3 = pp_28_56;
  assign pp_0_56_4 = pp_29_56;
  assign pp_0_56_5 = pp_30_56;
  assign pp_0_56_6 = pp_31_56;
  assign pp_0_57_0 = pp_26_57;
  assign pp_0_57_1 = pp_27_57;
  assign pp_0_57_2 = pp_28_57;
  assign pp_0_57_3 = pp_29_57;
  assign pp_0_57_4 = pp_30_57;
  assign pp_0_57_5 = pp_31_57;
  assign pp_0_58_0 = pp_27_58;
  assign pp_0_58_1 = pp_28_58;
  assign pp_0_58_2 = pp_29_58;
  assign pp_0_58_3 = pp_30_58;
  assign pp_0_58_4 = pp_31_58;
  assign pp_0_59_0 = pp_28_59;
  assign pp_0_59_1 = pp_29_59;
  assign pp_0_59_2 = pp_30_59;
  assign pp_0_59_3 = pp_31_59;
  assign pp_0_60_0 = pp_29_60;
  assign pp_0_60_1 = pp_30_60;
  assign pp_0_60_2 = pp_31_60;
  assign pp_0_61_0 = pp_30_61;
  assign pp_0_61_1 = pp_31_61;
  assign pp_0_62_0 = pp_31_62;

  assign pp_1_0_0 = pp_0_0_0;
  assign pp_1_1_0 = pp_0_1_0;
  assign pp_1_1_1 = pp_0_1_1;
  assign pp_1_2_0 = pp_0_2_0;
  assign pp_1_2_1 = pp_0_2_1;
  assign pp_1_2_2 = pp_0_2_2;
  assign pp_1_3_0 = pp_0_3_0;
  assign pp_1_3_1 = pp_0_3_1;
  assign pp_1_3_2 = pp_0_3_2;
  assign pp_1_3_3 = pp_0_3_3;
  MG_FA fa_0_4_0(
    .a(pp_0_4_0),
    .b(pp_0_4_1),
    .cin(pp_0_4_2),
    .sum(pp_1_4_0),
    .cout(pp_1_5_0)
  );

  assign pp_1_4_1 = pp_0_4_3;
  assign pp_1_4_2 = pp_0_4_4;
  assign pp_1_5_1 = pp_0_5_0;
  assign pp_1_5_2 = pp_0_5_1;
  assign pp_1_5_3 = pp_0_5_2;
  assign pp_1_5_4 = pp_0_5_3;
  assign pp_1_5_5 = pp_0_5_4;
  assign pp_1_5_6 = pp_0_5_5;
  MG_FA fa_0_6_0(
    .a(pp_0_6_0),
    .b(pp_0_6_1),
    .cin(pp_0_6_2),
    .sum(pp_1_6_0),
    .cout(pp_1_7_0)
  );

  assign pp_1_6_1 = pp_0_6_3;
  assign pp_1_6_2 = pp_0_6_4;
  assign pp_1_6_3 = pp_0_6_5;
  assign pp_1_6_4 = pp_0_6_6;
  MG_FA fa_0_7_0(
    .a(pp_0_7_0),
    .b(pp_0_7_1),
    .cin(pp_0_7_2),
    .sum(pp_1_7_1),
    .cout(pp_1_8_0)
  );

  MG_FA fa_0_7_1(
    .a(pp_0_7_3),
    .b(pp_0_7_4),
    .cin(pp_0_7_5),
    .sum(pp_1_7_2),
    .cout(pp_1_8_1)
  );

  assign pp_1_7_3 = pp_0_7_6;
  assign pp_1_7_4 = pp_0_7_7;
  assign pp_1_8_2 = pp_0_8_0;
  assign pp_1_8_3 = pp_0_8_1;
  assign pp_1_8_4 = pp_0_8_2;
  assign pp_1_8_5 = pp_0_8_3;
  assign pp_1_8_6 = pp_0_8_4;
  assign pp_1_8_7 = pp_0_8_5;
  assign pp_1_8_8 = pp_0_8_6;
  assign pp_1_8_9 = pp_0_8_7;
  assign pp_1_8_10 = pp_0_8_8;
  MG_FA fa_0_9_0(
    .a(pp_0_9_0),
    .b(pp_0_9_1),
    .cin(pp_0_9_2),
    .sum(pp_1_9_0),
    .cout(pp_1_10_0)
  );

  MG_FA fa_0_9_1(
    .a(pp_0_9_3),
    .b(pp_0_9_4),
    .cin(pp_0_9_5),
    .sum(pp_1_9_1),
    .cout(pp_1_10_1)
  );

  MG_HA ha_0_9_2(
    .a(pp_0_9_6),
    .b(pp_0_9_7),
    .sum(pp_1_9_2),
    .cout(pp_1_10_2)
  );

  assign pp_1_9_3 = pp_0_9_8;
  assign pp_1_9_4 = pp_0_9_9;
  MG_FA fa_0_10_0(
    .a(pp_0_10_0),
    .b(pp_0_10_1),
    .cin(pp_0_10_2),
    .sum(pp_1_10_3),
    .cout(pp_1_11_0)
  );

  MG_FA fa_0_10_1(
    .a(pp_0_10_3),
    .b(pp_0_10_4),
    .cin(pp_0_10_5),
    .sum(pp_1_10_4),
    .cout(pp_1_11_1)
  );

  MG_FA fa_0_10_2(
    .a(pp_0_10_6),
    .b(pp_0_10_7),
    .cin(pp_0_10_8),
    .sum(pp_1_10_5),
    .cout(pp_1_11_2)
  );

  assign pp_1_10_6 = pp_0_10_9;
  assign pp_1_10_7 = pp_0_10_10;
  MG_FA fa_0_11_0(
    .a(pp_0_11_0),
    .b(pp_0_11_1),
    .cin(pp_0_11_2),
    .sum(pp_1_11_3),
    .cout(pp_1_12_0)
  );

  MG_FA fa_0_11_1(
    .a(pp_0_11_3),
    .b(pp_0_11_4),
    .cin(pp_0_11_5),
    .sum(pp_1_11_4),
    .cout(pp_1_12_1)
  );

  MG_FA fa_0_11_2(
    .a(pp_0_11_6),
    .b(pp_0_11_7),
    .cin(pp_0_11_8),
    .sum(pp_1_11_5),
    .cout(pp_1_12_2)
  );

  MG_FA fa_0_11_3(
    .a(pp_0_11_9),
    .b(pp_0_11_10),
    .cin(pp_0_11_11),
    .sum(pp_1_11_6),
    .cout(pp_1_12_3)
  );

  MG_FA fa_0_12_0(
    .a(pp_0_12_0),
    .b(pp_0_12_1),
    .cin(pp_0_12_2),
    .sum(pp_1_12_4),
    .cout(pp_1_13_0)
  );

  MG_FA fa_0_12_1(
    .a(pp_0_12_3),
    .b(pp_0_12_4),
    .cin(pp_0_12_5),
    .sum(pp_1_12_5),
    .cout(pp_1_13_1)
  );

  MG_FA fa_0_12_2(
    .a(pp_0_12_6),
    .b(pp_0_12_7),
    .cin(pp_0_12_8),
    .sum(pp_1_12_6),
    .cout(pp_1_13_2)
  );

  MG_FA fa_0_12_3(
    .a(pp_0_12_9),
    .b(pp_0_12_10),
    .cin(pp_0_12_11),
    .sum(pp_1_12_7),
    .cout(pp_1_13_3)
  );

  assign pp_1_12_8 = pp_0_12_12;
  MG_FA fa_0_13_0(
    .a(pp_0_13_0),
    .b(pp_0_13_1),
    .cin(pp_0_13_2),
    .sum(pp_1_13_4),
    .cout(pp_1_14_0)
  );

  MG_FA fa_0_13_1(
    .a(pp_0_13_3),
    .b(pp_0_13_4),
    .cin(pp_0_13_5),
    .sum(pp_1_13_5),
    .cout(pp_1_14_1)
  );

  MG_FA fa_0_13_2(
    .a(pp_0_13_6),
    .b(pp_0_13_7),
    .cin(pp_0_13_8),
    .sum(pp_1_13_6),
    .cout(pp_1_14_2)
  );

  MG_FA fa_0_13_3(
    .a(pp_0_13_9),
    .b(pp_0_13_10),
    .cin(pp_0_13_11),
    .sum(pp_1_13_7),
    .cout(pp_1_14_3)
  );

  MG_HA ha_0_13_4(
    .a(pp_0_13_12),
    .b(pp_0_13_13),
    .sum(pp_1_13_8),
    .cout(pp_1_14_4)
  );

  MG_FA fa_0_14_0(
    .a(pp_0_14_0),
    .b(pp_0_14_1),
    .cin(pp_0_14_2),
    .sum(pp_1_14_5),
    .cout(pp_1_15_0)
  );

  MG_FA fa_0_14_1(
    .a(pp_0_14_3),
    .b(pp_0_14_4),
    .cin(pp_0_14_5),
    .sum(pp_1_14_6),
    .cout(pp_1_15_1)
  );

  MG_FA fa_0_14_2(
    .a(pp_0_14_6),
    .b(pp_0_14_7),
    .cin(pp_0_14_8),
    .sum(pp_1_14_7),
    .cout(pp_1_15_2)
  );

  MG_FA fa_0_14_3(
    .a(pp_0_14_9),
    .b(pp_0_14_10),
    .cin(pp_0_14_11),
    .sum(pp_1_14_8),
    .cout(pp_1_15_3)
  );

  MG_FA fa_0_14_4(
    .a(pp_0_14_12),
    .b(pp_0_14_13),
    .cin(pp_0_14_14),
    .sum(pp_1_14_9),
    .cout(pp_1_15_4)
  );

  MG_FA fa_0_15_0(
    .a(pp_0_15_0),
    .b(pp_0_15_1),
    .cin(pp_0_15_2),
    .sum(pp_1_15_5),
    .cout(pp_1_16_0)
  );

  MG_FA fa_0_15_1(
    .a(pp_0_15_3),
    .b(pp_0_15_4),
    .cin(pp_0_15_5),
    .sum(pp_1_15_6),
    .cout(pp_1_16_1)
  );

  MG_FA fa_0_15_2(
    .a(pp_0_15_6),
    .b(pp_0_15_7),
    .cin(pp_0_15_8),
    .sum(pp_1_15_7),
    .cout(pp_1_16_2)
  );

  MG_FA fa_0_15_3(
    .a(pp_0_15_9),
    .b(pp_0_15_10),
    .cin(pp_0_15_11),
    .sum(pp_1_15_8),
    .cout(pp_1_16_3)
  );

  MG_HA ha_0_15_4(
    .a(pp_0_15_12),
    .b(pp_0_15_13),
    .sum(pp_1_15_9),
    .cout(pp_1_16_4)
  );

  assign pp_1_15_10 = pp_0_15_14;
  assign pp_1_15_11 = pp_0_15_15;
  MG_FA fa_0_16_0(
    .a(pp_0_16_0),
    .b(pp_0_16_1),
    .cin(pp_0_16_2),
    .sum(pp_1_16_5),
    .cout(pp_1_17_0)
  );

  MG_FA fa_0_16_1(
    .a(pp_0_16_3),
    .b(pp_0_16_4),
    .cin(pp_0_16_5),
    .sum(pp_1_16_6),
    .cout(pp_1_17_1)
  );

  MG_FA fa_0_16_2(
    .a(pp_0_16_6),
    .b(pp_0_16_7),
    .cin(pp_0_16_8),
    .sum(pp_1_16_7),
    .cout(pp_1_17_2)
  );

  MG_FA fa_0_16_3(
    .a(pp_0_16_9),
    .b(pp_0_16_10),
    .cin(pp_0_16_11),
    .sum(pp_1_16_8),
    .cout(pp_1_17_3)
  );

  MG_FA fa_0_16_4(
    .a(pp_0_16_12),
    .b(pp_0_16_13),
    .cin(pp_0_16_14),
    .sum(pp_1_16_9),
    .cout(pp_1_17_4)
  );

  assign pp_1_16_10 = pp_0_16_15;
  assign pp_1_16_11 = pp_0_16_16;
  MG_FA fa_0_17_0(
    .a(pp_0_17_0),
    .b(pp_0_17_1),
    .cin(pp_0_17_2),
    .sum(pp_1_17_5),
    .cout(pp_1_18_0)
  );

  MG_FA fa_0_17_1(
    .a(pp_0_17_3),
    .b(pp_0_17_4),
    .cin(pp_0_17_5),
    .sum(pp_1_17_6),
    .cout(pp_1_18_1)
  );

  MG_FA fa_0_17_2(
    .a(pp_0_17_6),
    .b(pp_0_17_7),
    .cin(pp_0_17_8),
    .sum(pp_1_17_7),
    .cout(pp_1_18_2)
  );

  MG_FA fa_0_17_3(
    .a(pp_0_17_9),
    .b(pp_0_17_10),
    .cin(pp_0_17_11),
    .sum(pp_1_17_8),
    .cout(pp_1_18_3)
  );

  MG_FA fa_0_17_4(
    .a(pp_0_17_12),
    .b(pp_0_17_13),
    .cin(pp_0_17_14),
    .sum(pp_1_17_9),
    .cout(pp_1_18_4)
  );

  assign pp_1_17_10 = pp_0_17_15;
  assign pp_1_17_11 = pp_0_17_16;
  assign pp_1_17_12 = pp_0_17_17;
  MG_FA fa_0_18_0(
    .a(pp_0_18_0),
    .b(pp_0_18_1),
    .cin(pp_0_18_2),
    .sum(pp_1_18_5),
    .cout(pp_1_19_0)
  );

  MG_FA fa_0_18_1(
    .a(pp_0_18_3),
    .b(pp_0_18_4),
    .cin(pp_0_18_5),
    .sum(pp_1_18_6),
    .cout(pp_1_19_1)
  );

  MG_FA fa_0_18_2(
    .a(pp_0_18_6),
    .b(pp_0_18_7),
    .cin(pp_0_18_8),
    .sum(pp_1_18_7),
    .cout(pp_1_19_2)
  );

  MG_FA fa_0_18_3(
    .a(pp_0_18_9),
    .b(pp_0_18_10),
    .cin(pp_0_18_11),
    .sum(pp_1_18_8),
    .cout(pp_1_19_3)
  );

  MG_FA fa_0_18_4(
    .a(pp_0_18_12),
    .b(pp_0_18_13),
    .cin(pp_0_18_14),
    .sum(pp_1_18_9),
    .cout(pp_1_19_4)
  );

  MG_FA fa_0_18_5(
    .a(pp_0_18_15),
    .b(pp_0_18_16),
    .cin(pp_0_18_17),
    .sum(pp_1_18_10),
    .cout(pp_1_19_5)
  );

  assign pp_1_18_11 = pp_0_18_18;
  MG_FA fa_0_19_0(
    .a(pp_0_19_0),
    .b(pp_0_19_1),
    .cin(pp_0_19_2),
    .sum(pp_1_19_6),
    .cout(pp_1_20_0)
  );

  MG_FA fa_0_19_1(
    .a(pp_0_19_3),
    .b(pp_0_19_4),
    .cin(pp_0_19_5),
    .sum(pp_1_19_7),
    .cout(pp_1_20_1)
  );

  MG_FA fa_0_19_2(
    .a(pp_0_19_6),
    .b(pp_0_19_7),
    .cin(pp_0_19_8),
    .sum(pp_1_19_8),
    .cout(pp_1_20_2)
  );

  MG_FA fa_0_19_3(
    .a(pp_0_19_9),
    .b(pp_0_19_10),
    .cin(pp_0_19_11),
    .sum(pp_1_19_9),
    .cout(pp_1_20_3)
  );

  MG_FA fa_0_19_4(
    .a(pp_0_19_12),
    .b(pp_0_19_13),
    .cin(pp_0_19_14),
    .sum(pp_1_19_10),
    .cout(pp_1_20_4)
  );

  MG_FA fa_0_19_5(
    .a(pp_0_19_15),
    .b(pp_0_19_16),
    .cin(pp_0_19_17),
    .sum(pp_1_19_11),
    .cout(pp_1_20_5)
  );

  MG_HA ha_0_19_6(
    .a(pp_0_19_18),
    .b(pp_0_19_19),
    .sum(pp_1_19_12),
    .cout(pp_1_20_6)
  );

  MG_FA fa_0_20_0(
    .a(pp_0_20_0),
    .b(pp_0_20_1),
    .cin(pp_0_20_2),
    .sum(pp_1_20_7),
    .cout(pp_1_21_0)
  );

  MG_FA fa_0_20_1(
    .a(pp_0_20_3),
    .b(pp_0_20_4),
    .cin(pp_0_20_5),
    .sum(pp_1_20_8),
    .cout(pp_1_21_1)
  );

  MG_FA fa_0_20_2(
    .a(pp_0_20_6),
    .b(pp_0_20_7),
    .cin(pp_0_20_8),
    .sum(pp_1_20_9),
    .cout(pp_1_21_2)
  );

  MG_FA fa_0_20_3(
    .a(pp_0_20_9),
    .b(pp_0_20_10),
    .cin(pp_0_20_11),
    .sum(pp_1_20_10),
    .cout(pp_1_21_3)
  );

  MG_FA fa_0_20_4(
    .a(pp_0_20_12),
    .b(pp_0_20_13),
    .cin(pp_0_20_14),
    .sum(pp_1_20_11),
    .cout(pp_1_21_4)
  );

  MG_FA fa_0_20_5(
    .a(pp_0_20_15),
    .b(pp_0_20_16),
    .cin(pp_0_20_17),
    .sum(pp_1_20_12),
    .cout(pp_1_21_5)
  );

  MG_HA ha_0_20_6(
    .a(pp_0_20_18),
    .b(pp_0_20_19),
    .sum(pp_1_20_13),
    .cout(pp_1_21_6)
  );

  assign pp_1_20_14 = pp_0_20_20;
  MG_FA fa_0_21_0(
    .a(pp_0_21_0),
    .b(pp_0_21_1),
    .cin(pp_0_21_2),
    .sum(pp_1_21_7),
    .cout(pp_1_22_0)
  );

  MG_FA fa_0_21_1(
    .a(pp_0_21_3),
    .b(pp_0_21_4),
    .cin(pp_0_21_5),
    .sum(pp_1_21_8),
    .cout(pp_1_22_1)
  );

  MG_FA fa_0_21_2(
    .a(pp_0_21_6),
    .b(pp_0_21_7),
    .cin(pp_0_21_8),
    .sum(pp_1_21_9),
    .cout(pp_1_22_2)
  );

  MG_FA fa_0_21_3(
    .a(pp_0_21_9),
    .b(pp_0_21_10),
    .cin(pp_0_21_11),
    .sum(pp_1_21_10),
    .cout(pp_1_22_3)
  );

  MG_FA fa_0_21_4(
    .a(pp_0_21_12),
    .b(pp_0_21_13),
    .cin(pp_0_21_14),
    .sum(pp_1_21_11),
    .cout(pp_1_22_4)
  );

  MG_FA fa_0_21_5(
    .a(pp_0_21_15),
    .b(pp_0_21_16),
    .cin(pp_0_21_17),
    .sum(pp_1_21_12),
    .cout(pp_1_22_5)
  );

  MG_FA fa_0_21_6(
    .a(pp_0_21_18),
    .b(pp_0_21_19),
    .cin(pp_0_21_20),
    .sum(pp_1_21_13),
    .cout(pp_1_22_6)
  );

  assign pp_1_21_14 = pp_0_21_21;
  MG_FA fa_0_22_0(
    .a(pp_0_22_0),
    .b(pp_0_22_1),
    .cin(pp_0_22_2),
    .sum(pp_1_22_7),
    .cout(pp_1_23_0)
  );

  MG_FA fa_0_22_1(
    .a(pp_0_22_3),
    .b(pp_0_22_4),
    .cin(pp_0_22_5),
    .sum(pp_1_22_8),
    .cout(pp_1_23_1)
  );

  MG_FA fa_0_22_2(
    .a(pp_0_22_6),
    .b(pp_0_22_7),
    .cin(pp_0_22_8),
    .sum(pp_1_22_9),
    .cout(pp_1_23_2)
  );

  MG_FA fa_0_22_3(
    .a(pp_0_22_9),
    .b(pp_0_22_10),
    .cin(pp_0_22_11),
    .sum(pp_1_22_10),
    .cout(pp_1_23_3)
  );

  MG_FA fa_0_22_4(
    .a(pp_0_22_12),
    .b(pp_0_22_13),
    .cin(pp_0_22_14),
    .sum(pp_1_22_11),
    .cout(pp_1_23_4)
  );

  MG_FA fa_0_22_5(
    .a(pp_0_22_15),
    .b(pp_0_22_16),
    .cin(pp_0_22_17),
    .sum(pp_1_22_12),
    .cout(pp_1_23_5)
  );

  MG_FA fa_0_22_6(
    .a(pp_0_22_18),
    .b(pp_0_22_19),
    .cin(pp_0_22_20),
    .sum(pp_1_22_13),
    .cout(pp_1_23_6)
  );

  assign pp_1_22_14 = pp_0_22_21;
  assign pp_1_22_15 = pp_0_22_22;
  MG_FA fa_0_23_0(
    .a(pp_0_23_0),
    .b(pp_0_23_1),
    .cin(pp_0_23_2),
    .sum(pp_1_23_7),
    .cout(pp_1_24_0)
  );

  MG_FA fa_0_23_1(
    .a(pp_0_23_3),
    .b(pp_0_23_4),
    .cin(pp_0_23_5),
    .sum(pp_1_23_8),
    .cout(pp_1_24_1)
  );

  MG_FA fa_0_23_2(
    .a(pp_0_23_6),
    .b(pp_0_23_7),
    .cin(pp_0_23_8),
    .sum(pp_1_23_9),
    .cout(pp_1_24_2)
  );

  MG_FA fa_0_23_3(
    .a(pp_0_23_9),
    .b(pp_0_23_10),
    .cin(pp_0_23_11),
    .sum(pp_1_23_10),
    .cout(pp_1_24_3)
  );

  MG_FA fa_0_23_4(
    .a(pp_0_23_12),
    .b(pp_0_23_13),
    .cin(pp_0_23_14),
    .sum(pp_1_23_11),
    .cout(pp_1_24_4)
  );

  MG_FA fa_0_23_5(
    .a(pp_0_23_15),
    .b(pp_0_23_16),
    .cin(pp_0_23_17),
    .sum(pp_1_23_12),
    .cout(pp_1_24_5)
  );

  MG_FA fa_0_23_6(
    .a(pp_0_23_18),
    .b(pp_0_23_19),
    .cin(pp_0_23_20),
    .sum(pp_1_23_13),
    .cout(pp_1_24_6)
  );

  MG_FA fa_0_23_7(
    .a(pp_0_23_21),
    .b(pp_0_23_22),
    .cin(pp_0_23_23),
    .sum(pp_1_23_14),
    .cout(pp_1_24_7)
  );

  MG_FA fa_0_24_0(
    .a(pp_0_24_0),
    .b(pp_0_24_1),
    .cin(pp_0_24_2),
    .sum(pp_1_24_8),
    .cout(pp_1_25_0)
  );

  MG_FA fa_0_24_1(
    .a(pp_0_24_3),
    .b(pp_0_24_4),
    .cin(pp_0_24_5),
    .sum(pp_1_24_9),
    .cout(pp_1_25_1)
  );

  MG_FA fa_0_24_2(
    .a(pp_0_24_6),
    .b(pp_0_24_7),
    .cin(pp_0_24_8),
    .sum(pp_1_24_10),
    .cout(pp_1_25_2)
  );

  MG_FA fa_0_24_3(
    .a(pp_0_24_9),
    .b(pp_0_24_10),
    .cin(pp_0_24_11),
    .sum(pp_1_24_11),
    .cout(pp_1_25_3)
  );

  MG_FA fa_0_24_4(
    .a(pp_0_24_12),
    .b(pp_0_24_13),
    .cin(pp_0_24_14),
    .sum(pp_1_24_12),
    .cout(pp_1_25_4)
  );

  MG_FA fa_0_24_5(
    .a(pp_0_24_15),
    .b(pp_0_24_16),
    .cin(pp_0_24_17),
    .sum(pp_1_24_13),
    .cout(pp_1_25_5)
  );

  MG_FA fa_0_24_6(
    .a(pp_0_24_18),
    .b(pp_0_24_19),
    .cin(pp_0_24_20),
    .sum(pp_1_24_14),
    .cout(pp_1_25_6)
  );

  MG_FA fa_0_24_7(
    .a(pp_0_24_21),
    .b(pp_0_24_22),
    .cin(pp_0_24_23),
    .sum(pp_1_24_15),
    .cout(pp_1_25_7)
  );

  assign pp_1_24_16 = pp_0_24_24;
  assign pp_1_25_8 = pp_0_25_0;
  assign pp_1_25_9 = pp_0_25_1;
  assign pp_1_25_10 = pp_0_25_2;
  assign pp_1_25_11 = pp_0_25_3;
  assign pp_1_25_12 = pp_0_25_4;
  assign pp_1_25_13 = pp_0_25_5;
  assign pp_1_25_14 = pp_0_25_6;
  assign pp_1_25_15 = pp_0_25_7;
  assign pp_1_25_16 = pp_0_25_8;
  assign pp_1_25_17 = pp_0_25_9;
  assign pp_1_25_18 = pp_0_25_10;
  assign pp_1_25_19 = pp_0_25_11;
  assign pp_1_25_20 = pp_0_25_12;
  assign pp_1_25_21 = pp_0_25_13;
  assign pp_1_25_22 = pp_0_25_14;
  assign pp_1_25_23 = pp_0_25_15;
  assign pp_1_25_24 = pp_0_25_16;
  assign pp_1_25_25 = pp_0_25_17;
  assign pp_1_25_26 = pp_0_25_18;
  assign pp_1_25_27 = pp_0_25_19;
  assign pp_1_25_28 = pp_0_25_20;
  assign pp_1_25_29 = pp_0_25_21;
  assign pp_1_25_30 = pp_0_25_22;
  assign pp_1_25_31 = pp_0_25_23;
  assign pp_1_25_32 = pp_0_25_24;
  assign pp_1_25_33 = pp_0_25_25;
  MG_FA fa_0_26_0(
    .a(pp_0_26_0),
    .b(pp_0_26_1),
    .cin(pp_0_26_2),
    .sum(pp_1_26_0),
    .cout(pp_1_27_0)
  );

  MG_FA fa_0_26_1(
    .a(pp_0_26_3),
    .b(pp_0_26_4),
    .cin(pp_0_26_5),
    .sum(pp_1_26_1),
    .cout(pp_1_27_1)
  );

  MG_FA fa_0_26_2(
    .a(pp_0_26_6),
    .b(pp_0_26_7),
    .cin(pp_0_26_8),
    .sum(pp_1_26_2),
    .cout(pp_1_27_2)
  );

  MG_FA fa_0_26_3(
    .a(pp_0_26_9),
    .b(pp_0_26_10),
    .cin(pp_0_26_11),
    .sum(pp_1_26_3),
    .cout(pp_1_27_3)
  );

  MG_FA fa_0_26_4(
    .a(pp_0_26_12),
    .b(pp_0_26_13),
    .cin(pp_0_26_14),
    .sum(pp_1_26_4),
    .cout(pp_1_27_4)
  );

  MG_FA fa_0_26_5(
    .a(pp_0_26_15),
    .b(pp_0_26_16),
    .cin(pp_0_26_17),
    .sum(pp_1_26_5),
    .cout(pp_1_27_5)
  );

  MG_FA fa_0_26_6(
    .a(pp_0_26_18),
    .b(pp_0_26_19),
    .cin(pp_0_26_20),
    .sum(pp_1_26_6),
    .cout(pp_1_27_6)
  );

  MG_HA ha_0_26_7(
    .a(pp_0_26_21),
    .b(pp_0_26_22),
    .sum(pp_1_26_7),
    .cout(pp_1_27_7)
  );

  assign pp_1_26_8 = pp_0_26_23;
  assign pp_1_26_9 = pp_0_26_24;
  assign pp_1_26_10 = pp_0_26_25;
  assign pp_1_26_11 = pp_0_26_26;
  MG_FA fa_0_27_0(
    .a(pp_0_27_0),
    .b(pp_0_27_1),
    .cin(pp_0_27_2),
    .sum(pp_1_27_8),
    .cout(pp_1_28_0)
  );

  MG_FA fa_0_27_1(
    .a(pp_0_27_3),
    .b(pp_0_27_4),
    .cin(pp_0_27_5),
    .sum(pp_1_27_9),
    .cout(pp_1_28_1)
  );

  MG_FA fa_0_27_2(
    .a(pp_0_27_6),
    .b(pp_0_27_7),
    .cin(pp_0_27_8),
    .sum(pp_1_27_10),
    .cout(pp_1_28_2)
  );

  MG_FA fa_0_27_3(
    .a(pp_0_27_9),
    .b(pp_0_27_10),
    .cin(pp_0_27_11),
    .sum(pp_1_27_11),
    .cout(pp_1_28_3)
  );

  MG_FA fa_0_27_4(
    .a(pp_0_27_12),
    .b(pp_0_27_13),
    .cin(pp_0_27_14),
    .sum(pp_1_27_12),
    .cout(pp_1_28_4)
  );

  MG_FA fa_0_27_5(
    .a(pp_0_27_15),
    .b(pp_0_27_16),
    .cin(pp_0_27_17),
    .sum(pp_1_27_13),
    .cout(pp_1_28_5)
  );

  MG_FA fa_0_27_6(
    .a(pp_0_27_18),
    .b(pp_0_27_19),
    .cin(pp_0_27_20),
    .sum(pp_1_27_14),
    .cout(pp_1_28_6)
  );

  MG_FA fa_0_27_7(
    .a(pp_0_27_21),
    .b(pp_0_27_22),
    .cin(pp_0_27_23),
    .sum(pp_1_27_15),
    .cout(pp_1_28_7)
  );

  MG_FA fa_0_27_8(
    .a(pp_0_27_24),
    .b(pp_0_27_25),
    .cin(pp_0_27_26),
    .sum(pp_1_27_16),
    .cout(pp_1_28_8)
  );

  assign pp_1_27_17 = pp_0_27_27;
  MG_FA fa_0_28_0(
    .a(pp_0_28_0),
    .b(pp_0_28_1),
    .cin(pp_0_28_2),
    .sum(pp_1_28_9),
    .cout(pp_1_29_0)
  );

  MG_FA fa_0_28_1(
    .a(pp_0_28_3),
    .b(pp_0_28_4),
    .cin(pp_0_28_5),
    .sum(pp_1_28_10),
    .cout(pp_1_29_1)
  );

  MG_FA fa_0_28_2(
    .a(pp_0_28_6),
    .b(pp_0_28_7),
    .cin(pp_0_28_8),
    .sum(pp_1_28_11),
    .cout(pp_1_29_2)
  );

  MG_FA fa_0_28_3(
    .a(pp_0_28_9),
    .b(pp_0_28_10),
    .cin(pp_0_28_11),
    .sum(pp_1_28_12),
    .cout(pp_1_29_3)
  );

  MG_FA fa_0_28_4(
    .a(pp_0_28_12),
    .b(pp_0_28_13),
    .cin(pp_0_28_14),
    .sum(pp_1_28_13),
    .cout(pp_1_29_4)
  );

  MG_FA fa_0_28_5(
    .a(pp_0_28_15),
    .b(pp_0_28_16),
    .cin(pp_0_28_17),
    .sum(pp_1_28_14),
    .cout(pp_1_29_5)
  );

  MG_FA fa_0_28_6(
    .a(pp_0_28_18),
    .b(pp_0_28_19),
    .cin(pp_0_28_20),
    .sum(pp_1_28_15),
    .cout(pp_1_29_6)
  );

  MG_FA fa_0_28_7(
    .a(pp_0_28_21),
    .b(pp_0_28_22),
    .cin(pp_0_28_23),
    .sum(pp_1_28_16),
    .cout(pp_1_29_7)
  );

  MG_FA fa_0_28_8(
    .a(pp_0_28_24),
    .b(pp_0_28_25),
    .cin(pp_0_28_26),
    .sum(pp_1_28_17),
    .cout(pp_1_29_8)
  );

  assign pp_1_28_18 = pp_0_28_27;
  assign pp_1_28_19 = pp_0_28_28;
  MG_FA fa_0_29_0(
    .a(pp_0_29_0),
    .b(pp_0_29_1),
    .cin(pp_0_29_2),
    .sum(pp_1_29_9),
    .cout(pp_1_30_0)
  );

  MG_FA fa_0_29_1(
    .a(pp_0_29_3),
    .b(pp_0_29_4),
    .cin(pp_0_29_5),
    .sum(pp_1_29_10),
    .cout(pp_1_30_1)
  );

  MG_FA fa_0_29_2(
    .a(pp_0_29_6),
    .b(pp_0_29_7),
    .cin(pp_0_29_8),
    .sum(pp_1_29_11),
    .cout(pp_1_30_2)
  );

  MG_FA fa_0_29_3(
    .a(pp_0_29_9),
    .b(pp_0_29_10),
    .cin(pp_0_29_11),
    .sum(pp_1_29_12),
    .cout(pp_1_30_3)
  );

  MG_FA fa_0_29_4(
    .a(pp_0_29_12),
    .b(pp_0_29_13),
    .cin(pp_0_29_14),
    .sum(pp_1_29_13),
    .cout(pp_1_30_4)
  );

  MG_FA fa_0_29_5(
    .a(pp_0_29_15),
    .b(pp_0_29_16),
    .cin(pp_0_29_17),
    .sum(pp_1_29_14),
    .cout(pp_1_30_5)
  );

  MG_FA fa_0_29_6(
    .a(pp_0_29_18),
    .b(pp_0_29_19),
    .cin(pp_0_29_20),
    .sum(pp_1_29_15),
    .cout(pp_1_30_6)
  );

  MG_FA fa_0_29_7(
    .a(pp_0_29_21),
    .b(pp_0_29_22),
    .cin(pp_0_29_23),
    .sum(pp_1_29_16),
    .cout(pp_1_30_7)
  );

  MG_FA fa_0_29_8(
    .a(pp_0_29_24),
    .b(pp_0_29_25),
    .cin(pp_0_29_26),
    .sum(pp_1_29_17),
    .cout(pp_1_30_8)
  );

  MG_FA fa_0_29_9(
    .a(pp_0_29_27),
    .b(pp_0_29_28),
    .cin(pp_0_29_29),
    .sum(pp_1_29_18),
    .cout(pp_1_30_9)
  );

  MG_FA fa_0_30_0(
    .a(pp_0_30_0),
    .b(pp_0_30_1),
    .cin(pp_0_30_2),
    .sum(pp_1_30_10),
    .cout(pp_1_31_0)
  );

  MG_FA fa_0_30_1(
    .a(pp_0_30_3),
    .b(pp_0_30_4),
    .cin(pp_0_30_5),
    .sum(pp_1_30_11),
    .cout(pp_1_31_1)
  );

  MG_FA fa_0_30_2(
    .a(pp_0_30_6),
    .b(pp_0_30_7),
    .cin(pp_0_30_8),
    .sum(pp_1_30_12),
    .cout(pp_1_31_2)
  );

  MG_FA fa_0_30_3(
    .a(pp_0_30_9),
    .b(pp_0_30_10),
    .cin(pp_0_30_11),
    .sum(pp_1_30_13),
    .cout(pp_1_31_3)
  );

  MG_FA fa_0_30_4(
    .a(pp_0_30_12),
    .b(pp_0_30_13),
    .cin(pp_0_30_14),
    .sum(pp_1_30_14),
    .cout(pp_1_31_4)
  );

  MG_FA fa_0_30_5(
    .a(pp_0_30_15),
    .b(pp_0_30_16),
    .cin(pp_0_30_17),
    .sum(pp_1_30_15),
    .cout(pp_1_31_5)
  );

  MG_FA fa_0_30_6(
    .a(pp_0_30_18),
    .b(pp_0_30_19),
    .cin(pp_0_30_20),
    .sum(pp_1_30_16),
    .cout(pp_1_31_6)
  );

  MG_FA fa_0_30_7(
    .a(pp_0_30_21),
    .b(pp_0_30_22),
    .cin(pp_0_30_23),
    .sum(pp_1_30_17),
    .cout(pp_1_31_7)
  );

  MG_FA fa_0_30_8(
    .a(pp_0_30_24),
    .b(pp_0_30_25),
    .cin(pp_0_30_26),
    .sum(pp_1_30_18),
    .cout(pp_1_31_8)
  );

  MG_FA fa_0_30_9(
    .a(pp_0_30_27),
    .b(pp_0_30_28),
    .cin(pp_0_30_29),
    .sum(pp_1_30_19),
    .cout(pp_1_31_9)
  );

  assign pp_1_30_20 = pp_0_30_30;
  MG_FA fa_0_31_0(
    .a(pp_0_31_0),
    .b(pp_0_31_1),
    .cin(pp_0_31_2),
    .sum(pp_1_31_10),
    .cout(pp_1_32_0)
  );

  MG_FA fa_0_31_1(
    .a(pp_0_31_3),
    .b(pp_0_31_4),
    .cin(pp_0_31_5),
    .sum(pp_1_31_11),
    .cout(pp_1_32_1)
  );

  MG_FA fa_0_31_2(
    .a(pp_0_31_6),
    .b(pp_0_31_7),
    .cin(pp_0_31_8),
    .sum(pp_1_31_12),
    .cout(pp_1_32_2)
  );

  MG_FA fa_0_31_3(
    .a(pp_0_31_9),
    .b(pp_0_31_10),
    .cin(pp_0_31_11),
    .sum(pp_1_31_13),
    .cout(pp_1_32_3)
  );

  MG_FA fa_0_31_4(
    .a(pp_0_31_12),
    .b(pp_0_31_13),
    .cin(pp_0_31_14),
    .sum(pp_1_31_14),
    .cout(pp_1_32_4)
  );

  MG_FA fa_0_31_5(
    .a(pp_0_31_15),
    .b(pp_0_31_16),
    .cin(pp_0_31_17),
    .sum(pp_1_31_15),
    .cout(pp_1_32_5)
  );

  MG_FA fa_0_31_6(
    .a(pp_0_31_18),
    .b(pp_0_31_19),
    .cin(pp_0_31_20),
    .sum(pp_1_31_16),
    .cout(pp_1_32_6)
  );

  MG_FA fa_0_31_7(
    .a(pp_0_31_21),
    .b(pp_0_31_22),
    .cin(pp_0_31_23),
    .sum(pp_1_31_17),
    .cout(pp_1_32_7)
  );

  MG_FA fa_0_31_8(
    .a(pp_0_31_24),
    .b(pp_0_31_25),
    .cin(pp_0_31_26),
    .sum(pp_1_31_18),
    .cout(pp_1_32_8)
  );

  MG_FA fa_0_31_9(
    .a(pp_0_31_27),
    .b(pp_0_31_28),
    .cin(pp_0_31_29),
    .sum(pp_1_31_19),
    .cout(pp_1_32_9)
  );

  assign pp_1_31_20 = pp_0_31_30;
  assign pp_1_31_21 = pp_0_31_31;
  MG_FA fa_0_32_0(
    .a(pp_0_32_0),
    .b(pp_0_32_1),
    .cin(pp_0_32_2),
    .sum(pp_1_32_10),
    .cout(pp_1_33_0)
  );

  MG_FA fa_0_32_1(
    .a(pp_0_32_3),
    .b(pp_0_32_4),
    .cin(pp_0_32_5),
    .sum(pp_1_32_11),
    .cout(pp_1_33_1)
  );

  MG_FA fa_0_32_2(
    .a(pp_0_32_6),
    .b(pp_0_32_7),
    .cin(pp_0_32_8),
    .sum(pp_1_32_12),
    .cout(pp_1_33_2)
  );

  MG_FA fa_0_32_3(
    .a(pp_0_32_9),
    .b(pp_0_32_10),
    .cin(pp_0_32_11),
    .sum(pp_1_32_13),
    .cout(pp_1_33_3)
  );

  MG_FA fa_0_32_4(
    .a(pp_0_32_12),
    .b(pp_0_32_13),
    .cin(pp_0_32_14),
    .sum(pp_1_32_14),
    .cout(pp_1_33_4)
  );

  MG_FA fa_0_32_5(
    .a(pp_0_32_15),
    .b(pp_0_32_16),
    .cin(pp_0_32_17),
    .sum(pp_1_32_15),
    .cout(pp_1_33_5)
  );

  MG_FA fa_0_32_6(
    .a(pp_0_32_18),
    .b(pp_0_32_19),
    .cin(pp_0_32_20),
    .sum(pp_1_32_16),
    .cout(pp_1_33_6)
  );

  MG_FA fa_0_32_7(
    .a(pp_0_32_21),
    .b(pp_0_32_22),
    .cin(pp_0_32_23),
    .sum(pp_1_32_17),
    .cout(pp_1_33_7)
  );

  MG_FA fa_0_32_8(
    .a(pp_0_32_24),
    .b(pp_0_32_25),
    .cin(pp_0_32_26),
    .sum(pp_1_32_18),
    .cout(pp_1_33_8)
  );

  MG_FA fa_0_32_9(
    .a(pp_0_32_27),
    .b(pp_0_32_28),
    .cin(pp_0_32_29),
    .sum(pp_1_32_19),
    .cout(pp_1_33_9)
  );

  assign pp_1_32_20 = pp_0_32_30;
  MG_FA fa_0_33_0(
    .a(pp_0_33_0),
    .b(pp_0_33_1),
    .cin(pp_0_33_2),
    .sum(pp_1_33_10),
    .cout(pp_1_34_0)
  );

  MG_FA fa_0_33_1(
    .a(pp_0_33_3),
    .b(pp_0_33_4),
    .cin(pp_0_33_5),
    .sum(pp_1_33_11),
    .cout(pp_1_34_1)
  );

  MG_FA fa_0_33_2(
    .a(pp_0_33_6),
    .b(pp_0_33_7),
    .cin(pp_0_33_8),
    .sum(pp_1_33_12),
    .cout(pp_1_34_2)
  );

  MG_FA fa_0_33_3(
    .a(pp_0_33_9),
    .b(pp_0_33_10),
    .cin(pp_0_33_11),
    .sum(pp_1_33_13),
    .cout(pp_1_34_3)
  );

  MG_FA fa_0_33_4(
    .a(pp_0_33_12),
    .b(pp_0_33_13),
    .cin(pp_0_33_14),
    .sum(pp_1_33_14),
    .cout(pp_1_34_4)
  );

  MG_FA fa_0_33_5(
    .a(pp_0_33_15),
    .b(pp_0_33_16),
    .cin(pp_0_33_17),
    .sum(pp_1_33_15),
    .cout(pp_1_34_5)
  );

  MG_FA fa_0_33_6(
    .a(pp_0_33_18),
    .b(pp_0_33_19),
    .cin(pp_0_33_20),
    .sum(pp_1_33_16),
    .cout(pp_1_34_6)
  );

  MG_FA fa_0_33_7(
    .a(pp_0_33_21),
    .b(pp_0_33_22),
    .cin(pp_0_33_23),
    .sum(pp_1_33_17),
    .cout(pp_1_34_7)
  );

  MG_FA fa_0_33_8(
    .a(pp_0_33_24),
    .b(pp_0_33_25),
    .cin(pp_0_33_26),
    .sum(pp_1_33_18),
    .cout(pp_1_34_8)
  );

  MG_FA fa_0_33_9(
    .a(pp_0_33_27),
    .b(pp_0_33_28),
    .cin(pp_0_33_29),
    .sum(pp_1_33_19),
    .cout(pp_1_34_9)
  );

  MG_FA fa_0_34_0(
    .a(pp_0_34_0),
    .b(pp_0_34_1),
    .cin(pp_0_34_2),
    .sum(pp_1_34_10),
    .cout(pp_1_35_0)
  );

  MG_FA fa_0_34_1(
    .a(pp_0_34_3),
    .b(pp_0_34_4),
    .cin(pp_0_34_5),
    .sum(pp_1_34_11),
    .cout(pp_1_35_1)
  );

  MG_FA fa_0_34_2(
    .a(pp_0_34_6),
    .b(pp_0_34_7),
    .cin(pp_0_34_8),
    .sum(pp_1_34_12),
    .cout(pp_1_35_2)
  );

  MG_FA fa_0_34_3(
    .a(pp_0_34_9),
    .b(pp_0_34_10),
    .cin(pp_0_34_11),
    .sum(pp_1_34_13),
    .cout(pp_1_35_3)
  );

  MG_FA fa_0_34_4(
    .a(pp_0_34_12),
    .b(pp_0_34_13),
    .cin(pp_0_34_14),
    .sum(pp_1_34_14),
    .cout(pp_1_35_4)
  );

  MG_FA fa_0_34_5(
    .a(pp_0_34_15),
    .b(pp_0_34_16),
    .cin(pp_0_34_17),
    .sum(pp_1_34_15),
    .cout(pp_1_35_5)
  );

  MG_FA fa_0_34_6(
    .a(pp_0_34_18),
    .b(pp_0_34_19),
    .cin(pp_0_34_20),
    .sum(pp_1_34_16),
    .cout(pp_1_35_6)
  );

  MG_FA fa_0_34_7(
    .a(pp_0_34_21),
    .b(pp_0_34_22),
    .cin(pp_0_34_23),
    .sum(pp_1_34_17),
    .cout(pp_1_35_7)
  );

  MG_FA fa_0_34_8(
    .a(pp_0_34_24),
    .b(pp_0_34_25),
    .cin(pp_0_34_26),
    .sum(pp_1_34_18),
    .cout(pp_1_35_8)
  );

  assign pp_1_34_19 = pp_0_34_27;
  assign pp_1_34_20 = pp_0_34_28;
  MG_FA fa_0_35_0(
    .a(pp_0_35_0),
    .b(pp_0_35_1),
    .cin(pp_0_35_2),
    .sum(pp_1_35_9),
    .cout(pp_1_36_0)
  );

  MG_FA fa_0_35_1(
    .a(pp_0_35_3),
    .b(pp_0_35_4),
    .cin(pp_0_35_5),
    .sum(pp_1_35_10),
    .cout(pp_1_36_1)
  );

  MG_FA fa_0_35_2(
    .a(pp_0_35_6),
    .b(pp_0_35_7),
    .cin(pp_0_35_8),
    .sum(pp_1_35_11),
    .cout(pp_1_36_2)
  );

  MG_FA fa_0_35_3(
    .a(pp_0_35_9),
    .b(pp_0_35_10),
    .cin(pp_0_35_11),
    .sum(pp_1_35_12),
    .cout(pp_1_36_3)
  );

  MG_FA fa_0_35_4(
    .a(pp_0_35_12),
    .b(pp_0_35_13),
    .cin(pp_0_35_14),
    .sum(pp_1_35_13),
    .cout(pp_1_36_4)
  );

  MG_FA fa_0_35_5(
    .a(pp_0_35_15),
    .b(pp_0_35_16),
    .cin(pp_0_35_17),
    .sum(pp_1_35_14),
    .cout(pp_1_36_5)
  );

  MG_FA fa_0_35_6(
    .a(pp_0_35_18),
    .b(pp_0_35_19),
    .cin(pp_0_35_20),
    .sum(pp_1_35_15),
    .cout(pp_1_36_6)
  );

  MG_FA fa_0_35_7(
    .a(pp_0_35_21),
    .b(pp_0_35_22),
    .cin(pp_0_35_23),
    .sum(pp_1_35_16),
    .cout(pp_1_36_7)
  );

  MG_FA fa_0_35_8(
    .a(pp_0_35_24),
    .b(pp_0_35_25),
    .cin(pp_0_35_26),
    .sum(pp_1_35_17),
    .cout(pp_1_36_8)
  );

  assign pp_1_35_18 = pp_0_35_27;
  MG_FA fa_0_36_0(
    .a(pp_0_36_0),
    .b(pp_0_36_1),
    .cin(pp_0_36_2),
    .sum(pp_1_36_9),
    .cout(pp_1_37_0)
  );

  MG_FA fa_0_36_1(
    .a(pp_0_36_3),
    .b(pp_0_36_4),
    .cin(pp_0_36_5),
    .sum(pp_1_36_10),
    .cout(pp_1_37_1)
  );

  MG_FA fa_0_36_2(
    .a(pp_0_36_6),
    .b(pp_0_36_7),
    .cin(pp_0_36_8),
    .sum(pp_1_36_11),
    .cout(pp_1_37_2)
  );

  MG_FA fa_0_36_3(
    .a(pp_0_36_9),
    .b(pp_0_36_10),
    .cin(pp_0_36_11),
    .sum(pp_1_36_12),
    .cout(pp_1_37_3)
  );

  MG_FA fa_0_36_4(
    .a(pp_0_36_12),
    .b(pp_0_36_13),
    .cin(pp_0_36_14),
    .sum(pp_1_36_13),
    .cout(pp_1_37_4)
  );

  MG_FA fa_0_36_5(
    .a(pp_0_36_15),
    .b(pp_0_36_16),
    .cin(pp_0_36_17),
    .sum(pp_1_36_14),
    .cout(pp_1_37_5)
  );

  MG_FA fa_0_36_6(
    .a(pp_0_36_18),
    .b(pp_0_36_19),
    .cin(pp_0_36_20),
    .sum(pp_1_36_15),
    .cout(pp_1_37_6)
  );

  MG_FA fa_0_36_7(
    .a(pp_0_36_21),
    .b(pp_0_36_22),
    .cin(pp_0_36_23),
    .sum(pp_1_36_16),
    .cout(pp_1_37_7)
  );

  MG_FA fa_0_36_8(
    .a(pp_0_36_24),
    .b(pp_0_36_25),
    .cin(pp_0_36_26),
    .sum(pp_1_36_17),
    .cout(pp_1_37_8)
  );

  MG_FA fa_0_37_0(
    .a(pp_0_37_0),
    .b(pp_0_37_1),
    .cin(pp_0_37_2),
    .sum(pp_1_37_9),
    .cout(pp_1_38_0)
  );

  MG_FA fa_0_37_1(
    .a(pp_0_37_3),
    .b(pp_0_37_4),
    .cin(pp_0_37_5),
    .sum(pp_1_37_10),
    .cout(pp_1_38_1)
  );

  MG_FA fa_0_37_2(
    .a(pp_0_37_6),
    .b(pp_0_37_7),
    .cin(pp_0_37_8),
    .sum(pp_1_37_11),
    .cout(pp_1_38_2)
  );

  MG_FA fa_0_37_3(
    .a(pp_0_37_9),
    .b(pp_0_37_10),
    .cin(pp_0_37_11),
    .sum(pp_1_37_12),
    .cout(pp_1_38_3)
  );

  MG_FA fa_0_37_4(
    .a(pp_0_37_12),
    .b(pp_0_37_13),
    .cin(pp_0_37_14),
    .sum(pp_1_37_13),
    .cout(pp_1_38_4)
  );

  MG_FA fa_0_37_5(
    .a(pp_0_37_15),
    .b(pp_0_37_16),
    .cin(pp_0_37_17),
    .sum(pp_1_37_14),
    .cout(pp_1_38_5)
  );

  MG_FA fa_0_37_6(
    .a(pp_0_37_18),
    .b(pp_0_37_19),
    .cin(pp_0_37_20),
    .sum(pp_1_37_15),
    .cout(pp_1_38_6)
  );

  MG_FA fa_0_37_7(
    .a(pp_0_37_21),
    .b(pp_0_37_22),
    .cin(pp_0_37_23),
    .sum(pp_1_37_16),
    .cout(pp_1_38_7)
  );

  assign pp_1_37_17 = pp_0_37_24;
  assign pp_1_37_18 = pp_0_37_25;
  MG_FA fa_0_38_0(
    .a(pp_0_38_0),
    .b(pp_0_38_1),
    .cin(pp_0_38_2),
    .sum(pp_1_38_8),
    .cout(pp_1_39_0)
  );

  MG_FA fa_0_38_1(
    .a(pp_0_38_3),
    .b(pp_0_38_4),
    .cin(pp_0_38_5),
    .sum(pp_1_38_9),
    .cout(pp_1_39_1)
  );

  MG_FA fa_0_38_2(
    .a(pp_0_38_6),
    .b(pp_0_38_7),
    .cin(pp_0_38_8),
    .sum(pp_1_38_10),
    .cout(pp_1_39_2)
  );

  MG_FA fa_0_38_3(
    .a(pp_0_38_9),
    .b(pp_0_38_10),
    .cin(pp_0_38_11),
    .sum(pp_1_38_11),
    .cout(pp_1_39_3)
  );

  MG_FA fa_0_38_4(
    .a(pp_0_38_12),
    .b(pp_0_38_13),
    .cin(pp_0_38_14),
    .sum(pp_1_38_12),
    .cout(pp_1_39_4)
  );

  MG_FA fa_0_38_5(
    .a(pp_0_38_15),
    .b(pp_0_38_16),
    .cin(pp_0_38_17),
    .sum(pp_1_38_13),
    .cout(pp_1_39_5)
  );

  MG_FA fa_0_38_6(
    .a(pp_0_38_18),
    .b(pp_0_38_19),
    .cin(pp_0_38_20),
    .sum(pp_1_38_14),
    .cout(pp_1_39_6)
  );

  MG_FA fa_0_38_7(
    .a(pp_0_38_21),
    .b(pp_0_38_22),
    .cin(pp_0_38_23),
    .sum(pp_1_38_15),
    .cout(pp_1_39_7)
  );

  assign pp_1_38_16 = pp_0_38_24;
  MG_FA fa_0_39_0(
    .a(pp_0_39_0),
    .b(pp_0_39_1),
    .cin(pp_0_39_2),
    .sum(pp_1_39_8),
    .cout(pp_1_40_0)
  );

  MG_FA fa_0_39_1(
    .a(pp_0_39_3),
    .b(pp_0_39_4),
    .cin(pp_0_39_5),
    .sum(pp_1_39_9),
    .cout(pp_1_40_1)
  );

  MG_FA fa_0_39_2(
    .a(pp_0_39_6),
    .b(pp_0_39_7),
    .cin(pp_0_39_8),
    .sum(pp_1_39_10),
    .cout(pp_1_40_2)
  );

  MG_FA fa_0_39_3(
    .a(pp_0_39_9),
    .b(pp_0_39_10),
    .cin(pp_0_39_11),
    .sum(pp_1_39_11),
    .cout(pp_1_40_3)
  );

  MG_FA fa_0_39_4(
    .a(pp_0_39_12),
    .b(pp_0_39_13),
    .cin(pp_0_39_14),
    .sum(pp_1_39_12),
    .cout(pp_1_40_4)
  );

  MG_FA fa_0_39_5(
    .a(pp_0_39_15),
    .b(pp_0_39_16),
    .cin(pp_0_39_17),
    .sum(pp_1_39_13),
    .cout(pp_1_40_5)
  );

  MG_FA fa_0_39_6(
    .a(pp_0_39_18),
    .b(pp_0_39_19),
    .cin(pp_0_39_20),
    .sum(pp_1_39_14),
    .cout(pp_1_40_6)
  );

  MG_FA fa_0_39_7(
    .a(pp_0_39_21),
    .b(pp_0_39_22),
    .cin(pp_0_39_23),
    .sum(pp_1_39_15),
    .cout(pp_1_40_7)
  );

  MG_FA fa_0_40_0(
    .a(pp_0_40_0),
    .b(pp_0_40_1),
    .cin(pp_0_40_2),
    .sum(pp_1_40_8),
    .cout(pp_1_41_0)
  );

  MG_FA fa_0_40_1(
    .a(pp_0_40_3),
    .b(pp_0_40_4),
    .cin(pp_0_40_5),
    .sum(pp_1_40_9),
    .cout(pp_1_41_1)
  );

  MG_FA fa_0_40_2(
    .a(pp_0_40_6),
    .b(pp_0_40_7),
    .cin(pp_0_40_8),
    .sum(pp_1_40_10),
    .cout(pp_1_41_2)
  );

  MG_FA fa_0_40_3(
    .a(pp_0_40_9),
    .b(pp_0_40_10),
    .cin(pp_0_40_11),
    .sum(pp_1_40_11),
    .cout(pp_1_41_3)
  );

  MG_FA fa_0_40_4(
    .a(pp_0_40_12),
    .b(pp_0_40_13),
    .cin(pp_0_40_14),
    .sum(pp_1_40_12),
    .cout(pp_1_41_4)
  );

  assign pp_1_40_13 = pp_0_40_15;
  assign pp_1_40_14 = pp_0_40_16;
  assign pp_1_40_15 = pp_0_40_17;
  assign pp_1_40_16 = pp_0_40_18;
  assign pp_1_40_17 = pp_0_40_19;
  assign pp_1_40_18 = pp_0_40_20;
  assign pp_1_40_19 = pp_0_40_21;
  assign pp_1_40_20 = pp_0_40_22;
  MG_FA fa_0_41_0(
    .a(pp_0_41_0),
    .b(pp_0_41_1),
    .cin(pp_0_41_2),
    .sum(pp_1_41_5),
    .cout(pp_1_42_0)
  );

  MG_FA fa_0_41_1(
    .a(pp_0_41_3),
    .b(pp_0_41_4),
    .cin(pp_0_41_5),
    .sum(pp_1_41_6),
    .cout(pp_1_42_1)
  );

  MG_FA fa_0_41_2(
    .a(pp_0_41_6),
    .b(pp_0_41_7),
    .cin(pp_0_41_8),
    .sum(pp_1_41_7),
    .cout(pp_1_42_2)
  );

  MG_FA fa_0_41_3(
    .a(pp_0_41_9),
    .b(pp_0_41_10),
    .cin(pp_0_41_11),
    .sum(pp_1_41_8),
    .cout(pp_1_42_3)
  );

  MG_FA fa_0_41_4(
    .a(pp_0_41_12),
    .b(pp_0_41_13),
    .cin(pp_0_41_14),
    .sum(pp_1_41_9),
    .cout(pp_1_42_4)
  );

  MG_FA fa_0_41_5(
    .a(pp_0_41_15),
    .b(pp_0_41_16),
    .cin(pp_0_41_17),
    .sum(pp_1_41_10),
    .cout(pp_1_42_5)
  );

  assign pp_1_41_11 = pp_0_41_18;
  assign pp_1_41_12 = pp_0_41_19;
  assign pp_1_41_13 = pp_0_41_20;
  assign pp_1_41_14 = pp_0_41_21;
  MG_FA fa_0_42_0(
    .a(pp_0_42_0),
    .b(pp_0_42_1),
    .cin(pp_0_42_2),
    .sum(pp_1_42_6),
    .cout(pp_1_43_0)
  );

  MG_FA fa_0_42_1(
    .a(pp_0_42_3),
    .b(pp_0_42_4),
    .cin(pp_0_42_5),
    .sum(pp_1_42_7),
    .cout(pp_1_43_1)
  );

  MG_FA fa_0_42_2(
    .a(pp_0_42_6),
    .b(pp_0_42_7),
    .cin(pp_0_42_8),
    .sum(pp_1_42_8),
    .cout(pp_1_43_2)
  );

  MG_FA fa_0_42_3(
    .a(pp_0_42_9),
    .b(pp_0_42_10),
    .cin(pp_0_42_11),
    .sum(pp_1_42_9),
    .cout(pp_1_43_3)
  );

  MG_FA fa_0_42_4(
    .a(pp_0_42_12),
    .b(pp_0_42_13),
    .cin(pp_0_42_14),
    .sum(pp_1_42_10),
    .cout(pp_1_43_4)
  );

  MG_FA fa_0_42_5(
    .a(pp_0_42_15),
    .b(pp_0_42_16),
    .cin(pp_0_42_17),
    .sum(pp_1_42_11),
    .cout(pp_1_43_5)
  );

  MG_FA fa_0_42_6(
    .a(pp_0_42_18),
    .b(pp_0_42_19),
    .cin(pp_0_42_20),
    .sum(pp_1_42_12),
    .cout(pp_1_43_6)
  );

  MG_FA fa_0_43_0(
    .a(pp_0_43_0),
    .b(pp_0_43_1),
    .cin(pp_0_43_2),
    .sum(pp_1_43_7),
    .cout(pp_1_44_0)
  );

  MG_FA fa_0_43_1(
    .a(pp_0_43_3),
    .b(pp_0_43_4),
    .cin(pp_0_43_5),
    .sum(pp_1_43_8),
    .cout(pp_1_44_1)
  );

  MG_FA fa_0_43_2(
    .a(pp_0_43_6),
    .b(pp_0_43_7),
    .cin(pp_0_43_8),
    .sum(pp_1_43_9),
    .cout(pp_1_44_2)
  );

  MG_FA fa_0_43_3(
    .a(pp_0_43_9),
    .b(pp_0_43_10),
    .cin(pp_0_43_11),
    .sum(pp_1_43_10),
    .cout(pp_1_44_3)
  );

  MG_FA fa_0_43_4(
    .a(pp_0_43_12),
    .b(pp_0_43_13),
    .cin(pp_0_43_14),
    .sum(pp_1_43_11),
    .cout(pp_1_44_4)
  );

  MG_FA fa_0_43_5(
    .a(pp_0_43_15),
    .b(pp_0_43_16),
    .cin(pp_0_43_17),
    .sum(pp_1_43_12),
    .cout(pp_1_44_5)
  );

  assign pp_1_43_13 = pp_0_43_18;
  assign pp_1_43_14 = pp_0_43_19;
  assign pp_1_44_6 = pp_0_44_0;
  assign pp_1_44_7 = pp_0_44_1;
  assign pp_1_44_8 = pp_0_44_2;
  assign pp_1_44_9 = pp_0_44_3;
  assign pp_1_44_10 = pp_0_44_4;
  assign pp_1_44_11 = pp_0_44_5;
  assign pp_1_44_12 = pp_0_44_6;
  assign pp_1_44_13 = pp_0_44_7;
  assign pp_1_44_14 = pp_0_44_8;
  assign pp_1_44_15 = pp_0_44_9;
  assign pp_1_44_16 = pp_0_44_10;
  assign pp_1_44_17 = pp_0_44_11;
  assign pp_1_44_18 = pp_0_44_12;
  assign pp_1_44_19 = pp_0_44_13;
  assign pp_1_44_20 = pp_0_44_14;
  assign pp_1_44_21 = pp_0_44_15;
  assign pp_1_44_22 = pp_0_44_16;
  assign pp_1_44_23 = pp_0_44_17;
  assign pp_1_44_24 = pp_0_44_18;
  MG_FA fa_0_45_0(
    .a(pp_0_45_0),
    .b(pp_0_45_1),
    .cin(pp_0_45_2),
    .sum(pp_1_45_0),
    .cout(pp_1_46_0)
  );

  MG_FA fa_0_45_1(
    .a(pp_0_45_3),
    .b(pp_0_45_4),
    .cin(pp_0_45_5),
    .sum(pp_1_45_1),
    .cout(pp_1_46_1)
  );

  MG_FA fa_0_45_2(
    .a(pp_0_45_6),
    .b(pp_0_45_7),
    .cin(pp_0_45_8),
    .sum(pp_1_45_2),
    .cout(pp_1_46_2)
  );

  MG_FA fa_0_45_3(
    .a(pp_0_45_9),
    .b(pp_0_45_10),
    .cin(pp_0_45_11),
    .sum(pp_1_45_3),
    .cout(pp_1_46_3)
  );

  MG_FA fa_0_45_4(
    .a(pp_0_45_12),
    .b(pp_0_45_13),
    .cin(pp_0_45_14),
    .sum(pp_1_45_4),
    .cout(pp_1_46_4)
  );

  MG_FA fa_0_45_5(
    .a(pp_0_45_15),
    .b(pp_0_45_16),
    .cin(pp_0_45_17),
    .sum(pp_1_45_5),
    .cout(pp_1_46_5)
  );

  MG_FA fa_0_46_0(
    .a(pp_0_46_0),
    .b(pp_0_46_1),
    .cin(pp_0_46_2),
    .sum(pp_1_46_6),
    .cout(pp_1_47_0)
  );

  MG_FA fa_0_46_1(
    .a(pp_0_46_3),
    .b(pp_0_46_4),
    .cin(pp_0_46_5),
    .sum(pp_1_46_7),
    .cout(pp_1_47_1)
  );

  MG_FA fa_0_46_2(
    .a(pp_0_46_6),
    .b(pp_0_46_7),
    .cin(pp_0_46_8),
    .sum(pp_1_46_8),
    .cout(pp_1_47_2)
  );

  MG_FA fa_0_46_3(
    .a(pp_0_46_9),
    .b(pp_0_46_10),
    .cin(pp_0_46_11),
    .sum(pp_1_46_9),
    .cout(pp_1_47_3)
  );

  assign pp_1_46_10 = pp_0_46_12;
  assign pp_1_46_11 = pp_0_46_13;
  assign pp_1_46_12 = pp_0_46_14;
  assign pp_1_46_13 = pp_0_46_15;
  assign pp_1_46_14 = pp_0_46_16;
  MG_FA fa_0_47_0(
    .a(pp_0_47_0),
    .b(pp_0_47_1),
    .cin(pp_0_47_2),
    .sum(pp_1_47_4),
    .cout(pp_1_48_0)
  );

  MG_FA fa_0_47_1(
    .a(pp_0_47_3),
    .b(pp_0_47_4),
    .cin(pp_0_47_5),
    .sum(pp_1_47_5),
    .cout(pp_1_48_1)
  );

  MG_FA fa_0_47_2(
    .a(pp_0_47_6),
    .b(pp_0_47_7),
    .cin(pp_0_47_8),
    .sum(pp_1_47_6),
    .cout(pp_1_48_2)
  );

  MG_FA fa_0_47_3(
    .a(pp_0_47_9),
    .b(pp_0_47_10),
    .cin(pp_0_47_11),
    .sum(pp_1_47_7),
    .cout(pp_1_48_3)
  );

  assign pp_1_47_8 = pp_0_47_12;
  assign pp_1_47_9 = pp_0_47_13;
  assign pp_1_47_10 = pp_0_47_14;
  assign pp_1_47_11 = pp_0_47_15;
  MG_FA fa_0_48_0(
    .a(pp_0_48_0),
    .b(pp_0_48_1),
    .cin(pp_0_48_2),
    .sum(pp_1_48_4),
    .cout(pp_1_49_0)
  );

  MG_FA fa_0_48_1(
    .a(pp_0_48_3),
    .b(pp_0_48_4),
    .cin(pp_0_48_5),
    .sum(pp_1_48_5),
    .cout(pp_1_49_1)
  );

  MG_FA fa_0_48_2(
    .a(pp_0_48_6),
    .b(pp_0_48_7),
    .cin(pp_0_48_8),
    .sum(pp_1_48_6),
    .cout(pp_1_49_2)
  );

  MG_FA fa_0_48_3(
    .a(pp_0_48_9),
    .b(pp_0_48_10),
    .cin(pp_0_48_11),
    .sum(pp_1_48_7),
    .cout(pp_1_49_3)
  );

  MG_FA fa_0_48_4(
    .a(pp_0_48_12),
    .b(pp_0_48_13),
    .cin(pp_0_48_14),
    .sum(pp_1_48_8),
    .cout(pp_1_49_4)
  );

  MG_FA fa_0_49_0(
    .a(pp_0_49_0),
    .b(pp_0_49_1),
    .cin(pp_0_49_2),
    .sum(pp_1_49_5),
    .cout(pp_1_50_0)
  );

  MG_FA fa_0_49_1(
    .a(pp_0_49_3),
    .b(pp_0_49_4),
    .cin(pp_0_49_5),
    .sum(pp_1_49_6),
    .cout(pp_1_50_1)
  );

  MG_FA fa_0_49_2(
    .a(pp_0_49_6),
    .b(pp_0_49_7),
    .cin(pp_0_49_8),
    .sum(pp_1_49_7),
    .cout(pp_1_50_2)
  );

  MG_FA fa_0_49_3(
    .a(pp_0_49_9),
    .b(pp_0_49_10),
    .cin(pp_0_49_11),
    .sum(pp_1_49_8),
    .cout(pp_1_50_3)
  );

  assign pp_1_49_9 = pp_0_49_12;
  assign pp_1_49_10 = pp_0_49_13;
  MG_FA fa_0_50_0(
    .a(pp_0_50_0),
    .b(pp_0_50_1),
    .cin(pp_0_50_2),
    .sum(pp_1_50_4),
    .cout(pp_1_51_0)
  );

  MG_FA fa_0_50_1(
    .a(pp_0_50_3),
    .b(pp_0_50_4),
    .cin(pp_0_50_5),
    .sum(pp_1_50_5),
    .cout(pp_1_51_1)
  );

  MG_FA fa_0_50_2(
    .a(pp_0_50_6),
    .b(pp_0_50_7),
    .cin(pp_0_50_8),
    .sum(pp_1_50_6),
    .cout(pp_1_51_2)
  );

  MG_FA fa_0_50_3(
    .a(pp_0_50_9),
    .b(pp_0_50_10),
    .cin(pp_0_50_11),
    .sum(pp_1_50_7),
    .cout(pp_1_51_3)
  );

  assign pp_1_50_8 = pp_0_50_12;
  MG_FA fa_0_51_0(
    .a(pp_0_51_0),
    .b(pp_0_51_1),
    .cin(pp_0_51_2),
    .sum(pp_1_51_4),
    .cout(pp_1_52_0)
  );

  MG_FA fa_0_51_1(
    .a(pp_0_51_3),
    .b(pp_0_51_4),
    .cin(pp_0_51_5),
    .sum(pp_1_51_5),
    .cout(pp_1_52_1)
  );

  MG_FA fa_0_51_2(
    .a(pp_0_51_6),
    .b(pp_0_51_7),
    .cin(pp_0_51_8),
    .sum(pp_1_51_6),
    .cout(pp_1_52_2)
  );

  MG_FA fa_0_51_3(
    .a(pp_0_51_9),
    .b(pp_0_51_10),
    .cin(pp_0_51_11),
    .sum(pp_1_51_7),
    .cout(pp_1_52_3)
  );

  MG_FA fa_0_52_0(
    .a(pp_0_52_0),
    .b(pp_0_52_1),
    .cin(pp_0_52_2),
    .sum(pp_1_52_4),
    .cout(pp_1_53_0)
  );

  MG_FA fa_0_52_1(
    .a(pp_0_52_3),
    .b(pp_0_52_4),
    .cin(pp_0_52_5),
    .sum(pp_1_52_5),
    .cout(pp_1_53_1)
  );

  MG_FA fa_0_52_2(
    .a(pp_0_52_6),
    .b(pp_0_52_7),
    .cin(pp_0_52_8),
    .sum(pp_1_52_6),
    .cout(pp_1_53_2)
  );

  assign pp_1_52_7 = pp_0_52_9;
  assign pp_1_52_8 = pp_0_52_10;
  MG_FA fa_0_53_0(
    .a(pp_0_53_0),
    .b(pp_0_53_1),
    .cin(pp_0_53_2),
    .sum(pp_1_53_3),
    .cout(pp_1_54_0)
  );

  MG_FA fa_0_53_1(
    .a(pp_0_53_3),
    .b(pp_0_53_4),
    .cin(pp_0_53_5),
    .sum(pp_1_53_4),
    .cout(pp_1_54_1)
  );

  MG_FA fa_0_53_2(
    .a(pp_0_53_6),
    .b(pp_0_53_7),
    .cin(pp_0_53_8),
    .sum(pp_1_53_5),
    .cout(pp_1_54_2)
  );

  assign pp_1_53_6 = pp_0_53_9;
  MG_FA fa_0_54_0(
    .a(pp_0_54_0),
    .b(pp_0_54_1),
    .cin(pp_0_54_2),
    .sum(pp_1_54_3),
    .cout(pp_1_55_0)
  );

  MG_FA fa_0_54_1(
    .a(pp_0_54_3),
    .b(pp_0_54_4),
    .cin(pp_0_54_5),
    .sum(pp_1_54_4),
    .cout(pp_1_55_1)
  );

  MG_FA fa_0_54_2(
    .a(pp_0_54_6),
    .b(pp_0_54_7),
    .cin(pp_0_54_8),
    .sum(pp_1_54_5),
    .cout(pp_1_55_2)
  );

  MG_FA fa_0_55_0(
    .a(pp_0_55_0),
    .b(pp_0_55_1),
    .cin(pp_0_55_2),
    .sum(pp_1_55_3),
    .cout(pp_1_56_0)
  );

  MG_FA fa_0_55_1(
    .a(pp_0_55_3),
    .b(pp_0_55_4),
    .cin(pp_0_55_5),
    .sum(pp_1_55_4),
    .cout(pp_1_56_1)
  );

  assign pp_1_55_5 = pp_0_55_6;
  assign pp_1_55_6 = pp_0_55_7;
  assign pp_1_56_2 = pp_0_56_0;
  assign pp_1_56_3 = pp_0_56_1;
  assign pp_1_56_4 = pp_0_56_2;
  assign pp_1_56_5 = pp_0_56_3;
  assign pp_1_56_6 = pp_0_56_4;
  assign pp_1_56_7 = pp_0_56_5;
  assign pp_1_56_8 = pp_0_56_6;
  MG_FA fa_0_57_0(
    .a(pp_0_57_0),
    .b(pp_0_57_1),
    .cin(pp_0_57_2),
    .sum(pp_1_57_0),
    .cout(pp_1_58_0)
  );

  MG_FA fa_0_57_1(
    .a(pp_0_57_3),
    .b(pp_0_57_4),
    .cin(pp_0_57_5),
    .sum(pp_1_57_1),
    .cout(pp_1_58_1)
  );

  assign pp_1_58_2 = pp_0_58_0;
  assign pp_1_58_3 = pp_0_58_1;
  assign pp_1_58_4 = pp_0_58_2;
  assign pp_1_58_5 = pp_0_58_3;
  assign pp_1_58_6 = pp_0_58_4;
  assign pp_1_59_0 = pp_0_59_0;
  assign pp_1_59_1 = pp_0_59_1;
  assign pp_1_59_2 = pp_0_59_2;
  assign pp_1_59_3 = pp_0_59_3;
  MG_FA fa_0_60_0(
    .a(pp_0_60_0),
    .b(pp_0_60_1),
    .cin(pp_0_60_2),
    .sum(pp_1_60_0),
    .cout(pp_1_61_0)
  );

  assign pp_1_61_1 = pp_0_61_0;
  assign pp_1_61_2 = pp_0_61_1;
  assign pp_1_62_0 = pp_0_62_0;
  assign pp_2_0_0 = pp_1_0_0;
  assign pp_2_1_0 = pp_1_1_0;
  assign pp_2_1_1 = pp_1_1_1;
  assign pp_2_2_0 = pp_1_2_0;
  assign pp_2_2_1 = pp_1_2_1;
  assign pp_2_2_2 = pp_1_2_2;
  assign pp_2_3_0 = pp_1_3_0;
  assign pp_2_3_1 = pp_1_3_1;
  assign pp_2_3_2 = pp_1_3_2;
  assign pp_2_3_3 = pp_1_3_3;
  assign pp_2_4_0 = pp_1_4_0;
  assign pp_2_4_1 = pp_1_4_1;
  assign pp_2_4_2 = pp_1_4_2;
  MG_FA fa_1_5_0(
    .a(pp_1_5_0),
    .b(pp_1_5_1),
    .cin(pp_1_5_2),
    .sum(pp_2_5_0),
    .cout(pp_2_6_0)
  );

  MG_FA fa_1_5_1(
    .a(pp_1_5_3),
    .b(pp_1_5_4),
    .cin(pp_1_5_5),
    .sum(pp_2_5_1),
    .cout(pp_2_6_1)
  );

  assign pp_2_5_2 = pp_1_5_6;
  assign pp_2_6_2 = pp_1_6_0;
  assign pp_2_6_3 = pp_1_6_1;
  assign pp_2_6_4 = pp_1_6_2;
  assign pp_2_6_5 = pp_1_6_3;
  assign pp_2_6_6 = pp_1_6_4;
  MG_FA fa_1_7_0(
    .a(pp_1_7_0),
    .b(pp_1_7_1),
    .cin(pp_1_7_2),
    .sum(pp_2_7_0),
    .cout(pp_2_8_0)
  );

  MG_HA ha_1_7_1(
    .a(pp_1_7_3),
    .b(pp_1_7_4),
    .sum(pp_2_7_1),
    .cout(pp_2_8_1)
  );

  MG_FA fa_1_8_0(
    .a(pp_1_8_0),
    .b(pp_1_8_1),
    .cin(pp_1_8_2),
    .sum(pp_2_8_2),
    .cout(pp_2_9_0)
  );

  MG_FA fa_1_8_1(
    .a(pp_1_8_3),
    .b(pp_1_8_4),
    .cin(pp_1_8_5),
    .sum(pp_2_8_3),
    .cout(pp_2_9_1)
  );

  MG_FA fa_1_8_2(
    .a(pp_1_8_6),
    .b(pp_1_8_7),
    .cin(pp_1_8_8),
    .sum(pp_2_8_4),
    .cout(pp_2_9_2)
  );

  MG_HA ha_1_8_3(
    .a(pp_1_8_9),
    .b(pp_1_8_10),
    .sum(pp_2_8_5),
    .cout(pp_2_9_3)
  );

  assign pp_2_9_4 = pp_1_9_0;
  assign pp_2_9_5 = pp_1_9_1;
  assign pp_2_9_6 = pp_1_9_2;
  assign pp_2_9_7 = pp_1_9_3;
  assign pp_2_9_8 = pp_1_9_4;
  MG_FA fa_1_10_0(
    .a(pp_1_10_0),
    .b(pp_1_10_1),
    .cin(pp_1_10_2),
    .sum(pp_2_10_0),
    .cout(pp_2_11_0)
  );

  MG_FA fa_1_10_1(
    .a(pp_1_10_3),
    .b(pp_1_10_4),
    .cin(pp_1_10_5),
    .sum(pp_2_10_1),
    .cout(pp_2_11_1)
  );

  assign pp_2_10_2 = pp_1_10_6;
  assign pp_2_10_3 = pp_1_10_7;
  assign pp_2_11_2 = pp_1_11_0;
  assign pp_2_11_3 = pp_1_11_1;
  assign pp_2_11_4 = pp_1_11_2;
  assign pp_2_11_5 = pp_1_11_3;
  assign pp_2_11_6 = pp_1_11_4;
  assign pp_2_11_7 = pp_1_11_5;
  assign pp_2_11_8 = pp_1_11_6;
  MG_FA fa_1_12_0(
    .a(pp_1_12_0),
    .b(pp_1_12_1),
    .cin(pp_1_12_2),
    .sum(pp_2_12_0),
    .cout(pp_2_13_0)
  );

  MG_FA fa_1_12_1(
    .a(pp_1_12_3),
    .b(pp_1_12_4),
    .cin(pp_1_12_5),
    .sum(pp_2_12_1),
    .cout(pp_2_13_1)
  );

  MG_FA fa_1_12_2(
    .a(pp_1_12_6),
    .b(pp_1_12_7),
    .cin(pp_1_12_8),
    .sum(pp_2_12_2),
    .cout(pp_2_13_2)
  );

  MG_FA fa_1_13_0(
    .a(pp_1_13_0),
    .b(pp_1_13_1),
    .cin(pp_1_13_2),
    .sum(pp_2_13_3),
    .cout(pp_2_14_0)
  );

  MG_FA fa_1_13_1(
    .a(pp_1_13_3),
    .b(pp_1_13_4),
    .cin(pp_1_13_5),
    .sum(pp_2_13_4),
    .cout(pp_2_14_1)
  );

  MG_FA fa_1_13_2(
    .a(pp_1_13_6),
    .b(pp_1_13_7),
    .cin(pp_1_13_8),
    .sum(pp_2_13_5),
    .cout(pp_2_14_2)
  );

  assign pp_2_14_3 = pp_1_14_0;
  assign pp_2_14_4 = pp_1_14_1;
  assign pp_2_14_5 = pp_1_14_2;
  assign pp_2_14_6 = pp_1_14_3;
  assign pp_2_14_7 = pp_1_14_4;
  assign pp_2_14_8 = pp_1_14_5;
  assign pp_2_14_9 = pp_1_14_6;
  assign pp_2_14_10 = pp_1_14_7;
  assign pp_2_14_11 = pp_1_14_8;
  assign pp_2_14_12 = pp_1_14_9;
  MG_FA fa_1_15_0(
    .a(pp_1_15_0),
    .b(pp_1_15_1),
    .cin(pp_1_15_2),
    .sum(pp_2_15_0),
    .cout(pp_2_16_0)
  );

  MG_FA fa_1_15_1(
    .a(pp_1_15_3),
    .b(pp_1_15_4),
    .cin(pp_1_15_5),
    .sum(pp_2_15_1),
    .cout(pp_2_16_1)
  );

  MG_FA fa_1_15_2(
    .a(pp_1_15_6),
    .b(pp_1_15_7),
    .cin(pp_1_15_8),
    .sum(pp_2_15_2),
    .cout(pp_2_16_2)
  );

  MG_FA fa_1_15_3(
    .a(pp_1_15_9),
    .b(pp_1_15_10),
    .cin(pp_1_15_11),
    .sum(pp_2_15_3),
    .cout(pp_2_16_3)
  );

  MG_FA fa_1_16_0(
    .a(pp_1_16_0),
    .b(pp_1_16_1),
    .cin(pp_1_16_2),
    .sum(pp_2_16_4),
    .cout(pp_2_17_0)
  );

  MG_FA fa_1_16_1(
    .a(pp_1_16_3),
    .b(pp_1_16_4),
    .cin(pp_1_16_5),
    .sum(pp_2_16_5),
    .cout(pp_2_17_1)
  );

  MG_FA fa_1_16_2(
    .a(pp_1_16_6),
    .b(pp_1_16_7),
    .cin(pp_1_16_8),
    .sum(pp_2_16_6),
    .cout(pp_2_17_2)
  );

  MG_FA fa_1_16_3(
    .a(pp_1_16_9),
    .b(pp_1_16_10),
    .cin(pp_1_16_11),
    .sum(pp_2_16_7),
    .cout(pp_2_17_3)
  );

  MG_FA fa_1_17_0(
    .a(pp_1_17_0),
    .b(pp_1_17_1),
    .cin(pp_1_17_2),
    .sum(pp_2_17_4),
    .cout(pp_2_18_0)
  );

  MG_FA fa_1_17_1(
    .a(pp_1_17_3),
    .b(pp_1_17_4),
    .cin(pp_1_17_5),
    .sum(pp_2_17_5),
    .cout(pp_2_18_1)
  );

  MG_FA fa_1_17_2(
    .a(pp_1_17_6),
    .b(pp_1_17_7),
    .cin(pp_1_17_8),
    .sum(pp_2_17_6),
    .cout(pp_2_18_2)
  );

  MG_FA fa_1_17_3(
    .a(pp_1_17_9),
    .b(pp_1_17_10),
    .cin(pp_1_17_11),
    .sum(pp_2_17_7),
    .cout(pp_2_18_3)
  );

  assign pp_2_17_8 = pp_1_17_12;
  MG_FA fa_1_18_0(
    .a(pp_1_18_0),
    .b(pp_1_18_1),
    .cin(pp_1_18_2),
    .sum(pp_2_18_4),
    .cout(pp_2_19_0)
  );

  MG_FA fa_1_18_1(
    .a(pp_1_18_3),
    .b(pp_1_18_4),
    .cin(pp_1_18_5),
    .sum(pp_2_18_5),
    .cout(pp_2_19_1)
  );

  MG_FA fa_1_18_2(
    .a(pp_1_18_6),
    .b(pp_1_18_7),
    .cin(pp_1_18_8),
    .sum(pp_2_18_6),
    .cout(pp_2_19_2)
  );

  MG_FA fa_1_18_3(
    .a(pp_1_18_9),
    .b(pp_1_18_10),
    .cin(pp_1_18_11),
    .sum(pp_2_18_7),
    .cout(pp_2_19_3)
  );

  MG_FA fa_1_19_0(
    .a(pp_1_19_0),
    .b(pp_1_19_1),
    .cin(pp_1_19_2),
    .sum(pp_2_19_4),
    .cout(pp_2_20_0)
  );

  MG_FA fa_1_19_1(
    .a(pp_1_19_3),
    .b(pp_1_19_4),
    .cin(pp_1_19_5),
    .sum(pp_2_19_5),
    .cout(pp_2_20_1)
  );

  MG_FA fa_1_19_2(
    .a(pp_1_19_6),
    .b(pp_1_19_7),
    .cin(pp_1_19_8),
    .sum(pp_2_19_6),
    .cout(pp_2_20_2)
  );

  MG_FA fa_1_19_3(
    .a(pp_1_19_9),
    .b(pp_1_19_10),
    .cin(pp_1_19_11),
    .sum(pp_2_19_7),
    .cout(pp_2_20_3)
  );

  assign pp_2_19_8 = pp_1_19_12;
  MG_FA fa_1_20_0(
    .a(pp_1_20_0),
    .b(pp_1_20_1),
    .cin(pp_1_20_2),
    .sum(pp_2_20_4),
    .cout(pp_2_21_0)
  );

  MG_FA fa_1_20_1(
    .a(pp_1_20_3),
    .b(pp_1_20_4),
    .cin(pp_1_20_5),
    .sum(pp_2_20_5),
    .cout(pp_2_21_1)
  );

  MG_FA fa_1_20_2(
    .a(pp_1_20_6),
    .b(pp_1_20_7),
    .cin(pp_1_20_8),
    .sum(pp_2_20_6),
    .cout(pp_2_21_2)
  );

  MG_FA fa_1_20_3(
    .a(pp_1_20_9),
    .b(pp_1_20_10),
    .cin(pp_1_20_11),
    .sum(pp_2_20_7),
    .cout(pp_2_21_3)
  );

  MG_FA fa_1_20_4(
    .a(pp_1_20_12),
    .b(pp_1_20_13),
    .cin(pp_1_20_14),
    .sum(pp_2_20_8),
    .cout(pp_2_21_4)
  );

  MG_FA fa_1_21_0(
    .a(pp_1_21_0),
    .b(pp_1_21_1),
    .cin(pp_1_21_2),
    .sum(pp_2_21_5),
    .cout(pp_2_22_0)
  );

  MG_FA fa_1_21_1(
    .a(pp_1_21_3),
    .b(pp_1_21_4),
    .cin(pp_1_21_5),
    .sum(pp_2_21_6),
    .cout(pp_2_22_1)
  );

  MG_FA fa_1_21_2(
    .a(pp_1_21_6),
    .b(pp_1_21_7),
    .cin(pp_1_21_8),
    .sum(pp_2_21_7),
    .cout(pp_2_22_2)
  );

  MG_FA fa_1_21_3(
    .a(pp_1_21_9),
    .b(pp_1_21_10),
    .cin(pp_1_21_11),
    .sum(pp_2_21_8),
    .cout(pp_2_22_3)
  );

  MG_FA fa_1_21_4(
    .a(pp_1_21_12),
    .b(pp_1_21_13),
    .cin(pp_1_21_14),
    .sum(pp_2_21_9),
    .cout(pp_2_22_4)
  );

  assign pp_2_22_5 = pp_1_22_0;
  assign pp_2_22_6 = pp_1_22_1;
  assign pp_2_22_7 = pp_1_22_2;
  assign pp_2_22_8 = pp_1_22_3;
  assign pp_2_22_9 = pp_1_22_4;
  assign pp_2_22_10 = pp_1_22_5;
  assign pp_2_22_11 = pp_1_22_6;
  assign pp_2_22_12 = pp_1_22_7;
  assign pp_2_22_13 = pp_1_22_8;
  assign pp_2_22_14 = pp_1_22_9;
  assign pp_2_22_15 = pp_1_22_10;
  assign pp_2_22_16 = pp_1_22_11;
  assign pp_2_22_17 = pp_1_22_12;
  assign pp_2_22_18 = pp_1_22_13;
  assign pp_2_22_19 = pp_1_22_14;
  assign pp_2_22_20 = pp_1_22_15;
  MG_FA fa_1_23_0(
    .a(pp_1_23_0),
    .b(pp_1_23_1),
    .cin(pp_1_23_2),
    .sum(pp_2_23_0),
    .cout(pp_2_24_0)
  );

  MG_FA fa_1_23_1(
    .a(pp_1_23_3),
    .b(pp_1_23_4),
    .cin(pp_1_23_5),
    .sum(pp_2_23_1),
    .cout(pp_2_24_1)
  );

  MG_FA fa_1_23_2(
    .a(pp_1_23_6),
    .b(pp_1_23_7),
    .cin(pp_1_23_8),
    .sum(pp_2_23_2),
    .cout(pp_2_24_2)
  );

  MG_FA fa_1_23_3(
    .a(pp_1_23_9),
    .b(pp_1_23_10),
    .cin(pp_1_23_11),
    .sum(pp_2_23_3),
    .cout(pp_2_24_3)
  );

  MG_FA fa_1_23_4(
    .a(pp_1_23_12),
    .b(pp_1_23_13),
    .cin(pp_1_23_14),
    .sum(pp_2_23_4),
    .cout(pp_2_24_4)
  );

  MG_FA fa_1_24_0(
    .a(pp_1_24_0),
    .b(pp_1_24_1),
    .cin(pp_1_24_2),
    .sum(pp_2_24_5),
    .cout(pp_2_25_0)
  );

  MG_FA fa_1_24_1(
    .a(pp_1_24_3),
    .b(pp_1_24_4),
    .cin(pp_1_24_5),
    .sum(pp_2_24_6),
    .cout(pp_2_25_1)
  );

  MG_FA fa_1_24_2(
    .a(pp_1_24_6),
    .b(pp_1_24_7),
    .cin(pp_1_24_8),
    .sum(pp_2_24_7),
    .cout(pp_2_25_2)
  );

  MG_FA fa_1_24_3(
    .a(pp_1_24_9),
    .b(pp_1_24_10),
    .cin(pp_1_24_11),
    .sum(pp_2_24_8),
    .cout(pp_2_25_3)
  );

  MG_FA fa_1_24_4(
    .a(pp_1_24_12),
    .b(pp_1_24_13),
    .cin(pp_1_24_14),
    .sum(pp_2_24_9),
    .cout(pp_2_25_4)
  );

  assign pp_2_24_10 = pp_1_24_15;
  assign pp_2_24_11 = pp_1_24_16;
  MG_FA fa_1_25_0(
    .a(pp_1_25_0),
    .b(pp_1_25_1),
    .cin(pp_1_25_2),
    .sum(pp_2_25_5),
    .cout(pp_2_26_0)
  );

  MG_FA fa_1_25_1(
    .a(pp_1_25_3),
    .b(pp_1_25_4),
    .cin(pp_1_25_5),
    .sum(pp_2_25_6),
    .cout(pp_2_26_1)
  );

  MG_FA fa_1_25_2(
    .a(pp_1_25_6),
    .b(pp_1_25_7),
    .cin(pp_1_25_8),
    .sum(pp_2_25_7),
    .cout(pp_2_26_2)
  );

  MG_FA fa_1_25_3(
    .a(pp_1_25_9),
    .b(pp_1_25_10),
    .cin(pp_1_25_11),
    .sum(pp_2_25_8),
    .cout(pp_2_26_3)
  );

  MG_FA fa_1_25_4(
    .a(pp_1_25_12),
    .b(pp_1_25_13),
    .cin(pp_1_25_14),
    .sum(pp_2_25_9),
    .cout(pp_2_26_4)
  );

  MG_FA fa_1_25_5(
    .a(pp_1_25_15),
    .b(pp_1_25_16),
    .cin(pp_1_25_17),
    .sum(pp_2_25_10),
    .cout(pp_2_26_5)
  );

  MG_FA fa_1_25_6(
    .a(pp_1_25_18),
    .b(pp_1_25_19),
    .cin(pp_1_25_20),
    .sum(pp_2_25_11),
    .cout(pp_2_26_6)
  );

  MG_FA fa_1_25_7(
    .a(pp_1_25_21),
    .b(pp_1_25_22),
    .cin(pp_1_25_23),
    .sum(pp_2_25_12),
    .cout(pp_2_26_7)
  );

  MG_FA fa_1_25_8(
    .a(pp_1_25_24),
    .b(pp_1_25_25),
    .cin(pp_1_25_26),
    .sum(pp_2_25_13),
    .cout(pp_2_26_8)
  );

  MG_FA fa_1_25_9(
    .a(pp_1_25_27),
    .b(pp_1_25_28),
    .cin(pp_1_25_29),
    .sum(pp_2_25_14),
    .cout(pp_2_26_9)
  );

  MG_FA fa_1_25_10(
    .a(pp_1_25_30),
    .b(pp_1_25_31),
    .cin(pp_1_25_32),
    .sum(pp_2_25_15),
    .cout(pp_2_26_10)
  );

  assign pp_2_25_16 = pp_1_25_33;
  MG_FA fa_1_26_0(
    .a(pp_1_26_0),
    .b(pp_1_26_1),
    .cin(pp_1_26_2),
    .sum(pp_2_26_11),
    .cout(pp_2_27_0)
  );

  MG_FA fa_1_26_1(
    .a(pp_1_26_3),
    .b(pp_1_26_4),
    .cin(pp_1_26_5),
    .sum(pp_2_26_12),
    .cout(pp_2_27_1)
  );

  MG_FA fa_1_26_2(
    .a(pp_1_26_6),
    .b(pp_1_26_7),
    .cin(pp_1_26_8),
    .sum(pp_2_26_13),
    .cout(pp_2_27_2)
  );

  MG_FA fa_1_26_3(
    .a(pp_1_26_9),
    .b(pp_1_26_10),
    .cin(pp_1_26_11),
    .sum(pp_2_26_14),
    .cout(pp_2_27_3)
  );

  MG_FA fa_1_27_0(
    .a(pp_1_27_0),
    .b(pp_1_27_1),
    .cin(pp_1_27_2),
    .sum(pp_2_27_4),
    .cout(pp_2_28_0)
  );

  MG_FA fa_1_27_1(
    .a(pp_1_27_3),
    .b(pp_1_27_4),
    .cin(pp_1_27_5),
    .sum(pp_2_27_5),
    .cout(pp_2_28_1)
  );

  MG_FA fa_1_27_2(
    .a(pp_1_27_6),
    .b(pp_1_27_7),
    .cin(pp_1_27_8),
    .sum(pp_2_27_6),
    .cout(pp_2_28_2)
  );

  MG_FA fa_1_27_3(
    .a(pp_1_27_9),
    .b(pp_1_27_10),
    .cin(pp_1_27_11),
    .sum(pp_2_27_7),
    .cout(pp_2_28_3)
  );

  MG_FA fa_1_27_4(
    .a(pp_1_27_12),
    .b(pp_1_27_13),
    .cin(pp_1_27_14),
    .sum(pp_2_27_8),
    .cout(pp_2_28_4)
  );

  assign pp_2_27_9 = pp_1_27_15;
  assign pp_2_27_10 = pp_1_27_16;
  assign pp_2_27_11 = pp_1_27_17;
  MG_FA fa_1_28_0(
    .a(pp_1_28_0),
    .b(pp_1_28_1),
    .cin(pp_1_28_2),
    .sum(pp_2_28_5),
    .cout(pp_2_29_0)
  );

  MG_FA fa_1_28_1(
    .a(pp_1_28_3),
    .b(pp_1_28_4),
    .cin(pp_1_28_5),
    .sum(pp_2_28_6),
    .cout(pp_2_29_1)
  );

  MG_FA fa_1_28_2(
    .a(pp_1_28_6),
    .b(pp_1_28_7),
    .cin(pp_1_28_8),
    .sum(pp_2_28_7),
    .cout(pp_2_29_2)
  );

  MG_FA fa_1_28_3(
    .a(pp_1_28_9),
    .b(pp_1_28_10),
    .cin(pp_1_28_11),
    .sum(pp_2_28_8),
    .cout(pp_2_29_3)
  );

  MG_FA fa_1_28_4(
    .a(pp_1_28_12),
    .b(pp_1_28_13),
    .cin(pp_1_28_14),
    .sum(pp_2_28_9),
    .cout(pp_2_29_4)
  );

  MG_FA fa_1_28_5(
    .a(pp_1_28_15),
    .b(pp_1_28_16),
    .cin(pp_1_28_17),
    .sum(pp_2_28_10),
    .cout(pp_2_29_5)
  );

  assign pp_2_28_11 = pp_1_28_18;
  assign pp_2_28_12 = pp_1_28_19;
  MG_FA fa_1_29_0(
    .a(pp_1_29_0),
    .b(pp_1_29_1),
    .cin(pp_1_29_2),
    .sum(pp_2_29_6),
    .cout(pp_2_30_0)
  );

  MG_FA fa_1_29_1(
    .a(pp_1_29_3),
    .b(pp_1_29_4),
    .cin(pp_1_29_5),
    .sum(pp_2_29_7),
    .cout(pp_2_30_1)
  );

  MG_FA fa_1_29_2(
    .a(pp_1_29_6),
    .b(pp_1_29_7),
    .cin(pp_1_29_8),
    .sum(pp_2_29_8),
    .cout(pp_2_30_2)
  );

  MG_FA fa_1_29_3(
    .a(pp_1_29_9),
    .b(pp_1_29_10),
    .cin(pp_1_29_11),
    .sum(pp_2_29_9),
    .cout(pp_2_30_3)
  );

  MG_FA fa_1_29_4(
    .a(pp_1_29_12),
    .b(pp_1_29_13),
    .cin(pp_1_29_14),
    .sum(pp_2_29_10),
    .cout(pp_2_30_4)
  );

  MG_FA fa_1_29_5(
    .a(pp_1_29_15),
    .b(pp_1_29_16),
    .cin(pp_1_29_17),
    .sum(pp_2_29_11),
    .cout(pp_2_30_5)
  );

  assign pp_2_29_12 = pp_1_29_18;
  MG_FA fa_1_30_0(
    .a(pp_1_30_0),
    .b(pp_1_30_1),
    .cin(pp_1_30_2),
    .sum(pp_2_30_6),
    .cout(pp_2_31_0)
  );

  MG_FA fa_1_30_1(
    .a(pp_1_30_3),
    .b(pp_1_30_4),
    .cin(pp_1_30_5),
    .sum(pp_2_30_7),
    .cout(pp_2_31_1)
  );

  MG_FA fa_1_30_2(
    .a(pp_1_30_6),
    .b(pp_1_30_7),
    .cin(pp_1_30_8),
    .sum(pp_2_30_8),
    .cout(pp_2_31_2)
  );

  MG_FA fa_1_30_3(
    .a(pp_1_30_9),
    .b(pp_1_30_10),
    .cin(pp_1_30_11),
    .sum(pp_2_30_9),
    .cout(pp_2_31_3)
  );

  MG_FA fa_1_30_4(
    .a(pp_1_30_12),
    .b(pp_1_30_13),
    .cin(pp_1_30_14),
    .sum(pp_2_30_10),
    .cout(pp_2_31_4)
  );

  MG_FA fa_1_30_5(
    .a(pp_1_30_15),
    .b(pp_1_30_16),
    .cin(pp_1_30_17),
    .sum(pp_2_30_11),
    .cout(pp_2_31_5)
  );

  MG_FA fa_1_30_6(
    .a(pp_1_30_18),
    .b(pp_1_30_19),
    .cin(pp_1_30_20),
    .sum(pp_2_30_12),
    .cout(pp_2_31_6)
  );

  MG_FA fa_1_31_0(
    .a(pp_1_31_0),
    .b(pp_1_31_1),
    .cin(pp_1_31_2),
    .sum(pp_2_31_7),
    .cout(pp_2_32_0)
  );

  MG_FA fa_1_31_1(
    .a(pp_1_31_3),
    .b(pp_1_31_4),
    .cin(pp_1_31_5),
    .sum(pp_2_31_8),
    .cout(pp_2_32_1)
  );

  MG_FA fa_1_31_2(
    .a(pp_1_31_6),
    .b(pp_1_31_7),
    .cin(pp_1_31_8),
    .sum(pp_2_31_9),
    .cout(pp_2_32_2)
  );

  MG_FA fa_1_31_3(
    .a(pp_1_31_9),
    .b(pp_1_31_10),
    .cin(pp_1_31_11),
    .sum(pp_2_31_10),
    .cout(pp_2_32_3)
  );

  MG_FA fa_1_31_4(
    .a(pp_1_31_12),
    .b(pp_1_31_13),
    .cin(pp_1_31_14),
    .sum(pp_2_31_11),
    .cout(pp_2_32_4)
  );

  MG_FA fa_1_31_5(
    .a(pp_1_31_15),
    .b(pp_1_31_16),
    .cin(pp_1_31_17),
    .sum(pp_2_31_12),
    .cout(pp_2_32_5)
  );

  MG_FA fa_1_31_6(
    .a(pp_1_31_18),
    .b(pp_1_31_19),
    .cin(pp_1_31_20),
    .sum(pp_2_31_13),
    .cout(pp_2_32_6)
  );

  assign pp_2_31_14 = pp_1_31_21;
  MG_FA fa_1_32_0(
    .a(pp_1_32_0),
    .b(pp_1_32_1),
    .cin(pp_1_32_2),
    .sum(pp_2_32_7),
    .cout(pp_2_33_0)
  );

  MG_FA fa_1_32_1(
    .a(pp_1_32_3),
    .b(pp_1_32_4),
    .cin(pp_1_32_5),
    .sum(pp_2_32_8),
    .cout(pp_2_33_1)
  );

  MG_FA fa_1_32_2(
    .a(pp_1_32_6),
    .b(pp_1_32_7),
    .cin(pp_1_32_8),
    .sum(pp_2_32_9),
    .cout(pp_2_33_2)
  );

  MG_FA fa_1_32_3(
    .a(pp_1_32_9),
    .b(pp_1_32_10),
    .cin(pp_1_32_11),
    .sum(pp_2_32_10),
    .cout(pp_2_33_3)
  );

  MG_FA fa_1_32_4(
    .a(pp_1_32_12),
    .b(pp_1_32_13),
    .cin(pp_1_32_14),
    .sum(pp_2_32_11),
    .cout(pp_2_33_4)
  );

  MG_FA fa_1_32_5(
    .a(pp_1_32_15),
    .b(pp_1_32_16),
    .cin(pp_1_32_17),
    .sum(pp_2_32_12),
    .cout(pp_2_33_5)
  );

  MG_FA fa_1_32_6(
    .a(pp_1_32_18),
    .b(pp_1_32_19),
    .cin(pp_1_32_20),
    .sum(pp_2_32_13),
    .cout(pp_2_33_6)
  );

  MG_FA fa_1_33_0(
    .a(pp_1_33_0),
    .b(pp_1_33_1),
    .cin(pp_1_33_2),
    .sum(pp_2_33_7),
    .cout(pp_2_34_0)
  );

  MG_FA fa_1_33_1(
    .a(pp_1_33_3),
    .b(pp_1_33_4),
    .cin(pp_1_33_5),
    .sum(pp_2_33_8),
    .cout(pp_2_34_1)
  );

  MG_FA fa_1_33_2(
    .a(pp_1_33_6),
    .b(pp_1_33_7),
    .cin(pp_1_33_8),
    .sum(pp_2_33_9),
    .cout(pp_2_34_2)
  );

  MG_FA fa_1_33_3(
    .a(pp_1_33_9),
    .b(pp_1_33_10),
    .cin(pp_1_33_11),
    .sum(pp_2_33_10),
    .cout(pp_2_34_3)
  );

  MG_FA fa_1_33_4(
    .a(pp_1_33_12),
    .b(pp_1_33_13),
    .cin(pp_1_33_14),
    .sum(pp_2_33_11),
    .cout(pp_2_34_4)
  );

  MG_FA fa_1_33_5(
    .a(pp_1_33_15),
    .b(pp_1_33_16),
    .cin(pp_1_33_17),
    .sum(pp_2_33_12),
    .cout(pp_2_34_5)
  );

  assign pp_2_33_13 = pp_1_33_18;
  assign pp_2_33_14 = pp_1_33_19;
  MG_FA fa_1_34_0(
    .a(pp_1_34_0),
    .b(pp_1_34_1),
    .cin(pp_1_34_2),
    .sum(pp_2_34_6),
    .cout(pp_2_35_0)
  );

  MG_FA fa_1_34_1(
    .a(pp_1_34_3),
    .b(pp_1_34_4),
    .cin(pp_1_34_5),
    .sum(pp_2_34_7),
    .cout(pp_2_35_1)
  );

  MG_FA fa_1_34_2(
    .a(pp_1_34_6),
    .b(pp_1_34_7),
    .cin(pp_1_34_8),
    .sum(pp_2_34_8),
    .cout(pp_2_35_2)
  );

  MG_FA fa_1_34_3(
    .a(pp_1_34_9),
    .b(pp_1_34_10),
    .cin(pp_1_34_11),
    .sum(pp_2_34_9),
    .cout(pp_2_35_3)
  );

  MG_FA fa_1_34_4(
    .a(pp_1_34_12),
    .b(pp_1_34_13),
    .cin(pp_1_34_14),
    .sum(pp_2_34_10),
    .cout(pp_2_35_4)
  );

  MG_FA fa_1_34_5(
    .a(pp_1_34_15),
    .b(pp_1_34_16),
    .cin(pp_1_34_17),
    .sum(pp_2_34_11),
    .cout(pp_2_35_5)
  );

  MG_FA fa_1_34_6(
    .a(pp_1_34_18),
    .b(pp_1_34_19),
    .cin(pp_1_34_20),
    .sum(pp_2_34_12),
    .cout(pp_2_35_6)
  );

  MG_FA fa_1_35_0(
    .a(pp_1_35_0),
    .b(pp_1_35_1),
    .cin(pp_1_35_2),
    .sum(pp_2_35_7),
    .cout(pp_2_36_0)
  );

  MG_FA fa_1_35_1(
    .a(pp_1_35_3),
    .b(pp_1_35_4),
    .cin(pp_1_35_5),
    .sum(pp_2_35_8),
    .cout(pp_2_36_1)
  );

  MG_FA fa_1_35_2(
    .a(pp_1_35_6),
    .b(pp_1_35_7),
    .cin(pp_1_35_8),
    .sum(pp_2_35_9),
    .cout(pp_2_36_2)
  );

  MG_FA fa_1_35_3(
    .a(pp_1_35_9),
    .b(pp_1_35_10),
    .cin(pp_1_35_11),
    .sum(pp_2_35_10),
    .cout(pp_2_36_3)
  );

  MG_FA fa_1_35_4(
    .a(pp_1_35_12),
    .b(pp_1_35_13),
    .cin(pp_1_35_14),
    .sum(pp_2_35_11),
    .cout(pp_2_36_4)
  );

  MG_FA fa_1_35_5(
    .a(pp_1_35_15),
    .b(pp_1_35_16),
    .cin(pp_1_35_17),
    .sum(pp_2_35_12),
    .cout(pp_2_36_5)
  );

  assign pp_2_35_13 = pp_1_35_18;
  MG_FA fa_1_36_0(
    .a(pp_1_36_0),
    .b(pp_1_36_1),
    .cin(pp_1_36_2),
    .sum(pp_2_36_6),
    .cout(pp_2_37_0)
  );

  MG_FA fa_1_36_1(
    .a(pp_1_36_3),
    .b(pp_1_36_4),
    .cin(pp_1_36_5),
    .sum(pp_2_36_7),
    .cout(pp_2_37_1)
  );

  MG_FA fa_1_36_2(
    .a(pp_1_36_6),
    .b(pp_1_36_7),
    .cin(pp_1_36_8),
    .sum(pp_2_36_8),
    .cout(pp_2_37_2)
  );

  MG_FA fa_1_36_3(
    .a(pp_1_36_9),
    .b(pp_1_36_10),
    .cin(pp_1_36_11),
    .sum(pp_2_36_9),
    .cout(pp_2_37_3)
  );

  MG_FA fa_1_36_4(
    .a(pp_1_36_12),
    .b(pp_1_36_13),
    .cin(pp_1_36_14),
    .sum(pp_2_36_10),
    .cout(pp_2_37_4)
  );

  MG_FA fa_1_36_5(
    .a(pp_1_36_15),
    .b(pp_1_36_16),
    .cin(pp_1_36_17),
    .sum(pp_2_36_11),
    .cout(pp_2_37_5)
  );

  MG_FA fa_1_37_0(
    .a(pp_1_37_0),
    .b(pp_1_37_1),
    .cin(pp_1_37_2),
    .sum(pp_2_37_6),
    .cout(pp_2_38_0)
  );

  MG_FA fa_1_37_1(
    .a(pp_1_37_3),
    .b(pp_1_37_4),
    .cin(pp_1_37_5),
    .sum(pp_2_37_7),
    .cout(pp_2_38_1)
  );

  MG_FA fa_1_37_2(
    .a(pp_1_37_6),
    .b(pp_1_37_7),
    .cin(pp_1_37_8),
    .sum(pp_2_37_8),
    .cout(pp_2_38_2)
  );

  MG_FA fa_1_37_3(
    .a(pp_1_37_9),
    .b(pp_1_37_10),
    .cin(pp_1_37_11),
    .sum(pp_2_37_9),
    .cout(pp_2_38_3)
  );

  MG_FA fa_1_37_4(
    .a(pp_1_37_12),
    .b(pp_1_37_13),
    .cin(pp_1_37_14),
    .sum(pp_2_37_10),
    .cout(pp_2_38_4)
  );

  MG_FA fa_1_37_5(
    .a(pp_1_37_15),
    .b(pp_1_37_16),
    .cin(pp_1_37_17),
    .sum(pp_2_37_11),
    .cout(pp_2_38_5)
  );

  assign pp_2_37_12 = pp_1_37_18;
  MG_FA fa_1_38_0(
    .a(pp_1_38_0),
    .b(pp_1_38_1),
    .cin(pp_1_38_2),
    .sum(pp_2_38_6),
    .cout(pp_2_39_0)
  );

  MG_FA fa_1_38_1(
    .a(pp_1_38_3),
    .b(pp_1_38_4),
    .cin(pp_1_38_5),
    .sum(pp_2_38_7),
    .cout(pp_2_39_1)
  );

  MG_FA fa_1_38_2(
    .a(pp_1_38_6),
    .b(pp_1_38_7),
    .cin(pp_1_38_8),
    .sum(pp_2_38_8),
    .cout(pp_2_39_2)
  );

  MG_FA fa_1_38_3(
    .a(pp_1_38_9),
    .b(pp_1_38_10),
    .cin(pp_1_38_11),
    .sum(pp_2_38_9),
    .cout(pp_2_39_3)
  );

  MG_FA fa_1_38_4(
    .a(pp_1_38_12),
    .b(pp_1_38_13),
    .cin(pp_1_38_14),
    .sum(pp_2_38_10),
    .cout(pp_2_39_4)
  );

  assign pp_2_38_11 = pp_1_38_15;
  assign pp_2_38_12 = pp_1_38_16;
  MG_FA fa_1_39_0(
    .a(pp_1_39_0),
    .b(pp_1_39_1),
    .cin(pp_1_39_2),
    .sum(pp_2_39_5),
    .cout(pp_2_40_0)
  );

  MG_FA fa_1_39_1(
    .a(pp_1_39_3),
    .b(pp_1_39_4),
    .cin(pp_1_39_5),
    .sum(pp_2_39_6),
    .cout(pp_2_40_1)
  );

  MG_FA fa_1_39_2(
    .a(pp_1_39_6),
    .b(pp_1_39_7),
    .cin(pp_1_39_8),
    .sum(pp_2_39_7),
    .cout(pp_2_40_2)
  );

  MG_FA fa_1_39_3(
    .a(pp_1_39_9),
    .b(pp_1_39_10),
    .cin(pp_1_39_11),
    .sum(pp_2_39_8),
    .cout(pp_2_40_3)
  );

  MG_FA fa_1_39_4(
    .a(pp_1_39_12),
    .b(pp_1_39_13),
    .cin(pp_1_39_14),
    .sum(pp_2_39_9),
    .cout(pp_2_40_4)
  );

  assign pp_2_39_10 = pp_1_39_15;
  MG_FA fa_1_40_0(
    .a(pp_1_40_0),
    .b(pp_1_40_1),
    .cin(pp_1_40_2),
    .sum(pp_2_40_5),
    .cout(pp_2_41_0)
  );

  MG_FA fa_1_40_1(
    .a(pp_1_40_3),
    .b(pp_1_40_4),
    .cin(pp_1_40_5),
    .sum(pp_2_40_6),
    .cout(pp_2_41_1)
  );

  MG_FA fa_1_40_2(
    .a(pp_1_40_6),
    .b(pp_1_40_7),
    .cin(pp_1_40_8),
    .sum(pp_2_40_7),
    .cout(pp_2_41_2)
  );

  MG_FA fa_1_40_3(
    .a(pp_1_40_9),
    .b(pp_1_40_10),
    .cin(pp_1_40_11),
    .sum(pp_2_40_8),
    .cout(pp_2_41_3)
  );

  MG_FA fa_1_40_4(
    .a(pp_1_40_12),
    .b(pp_1_40_13),
    .cin(pp_1_40_14),
    .sum(pp_2_40_9),
    .cout(pp_2_41_4)
  );

  MG_FA fa_1_40_5(
    .a(pp_1_40_15),
    .b(pp_1_40_16),
    .cin(pp_1_40_17),
    .sum(pp_2_40_10),
    .cout(pp_2_41_5)
  );

  MG_FA fa_1_40_6(
    .a(pp_1_40_18),
    .b(pp_1_40_19),
    .cin(pp_1_40_20),
    .sum(pp_2_40_11),
    .cout(pp_2_41_6)
  );

  MG_FA fa_1_41_0(
    .a(pp_1_41_0),
    .b(pp_1_41_1),
    .cin(pp_1_41_2),
    .sum(pp_2_41_7),
    .cout(pp_2_42_0)
  );

  MG_FA fa_1_41_1(
    .a(pp_1_41_3),
    .b(pp_1_41_4),
    .cin(pp_1_41_5),
    .sum(pp_2_41_8),
    .cout(pp_2_42_1)
  );

  MG_FA fa_1_41_2(
    .a(pp_1_41_6),
    .b(pp_1_41_7),
    .cin(pp_1_41_8),
    .sum(pp_2_41_9),
    .cout(pp_2_42_2)
  );

  MG_FA fa_1_41_3(
    .a(pp_1_41_9),
    .b(pp_1_41_10),
    .cin(pp_1_41_11),
    .sum(pp_2_41_10),
    .cout(pp_2_42_3)
  );

  MG_FA fa_1_41_4(
    .a(pp_1_41_12),
    .b(pp_1_41_13),
    .cin(pp_1_41_14),
    .sum(pp_2_41_11),
    .cout(pp_2_42_4)
  );

  MG_FA fa_1_42_0(
    .a(pp_1_42_0),
    .b(pp_1_42_1),
    .cin(pp_1_42_2),
    .sum(pp_2_42_5),
    .cout(pp_2_43_0)
  );

  MG_FA fa_1_42_1(
    .a(pp_1_42_3),
    .b(pp_1_42_4),
    .cin(pp_1_42_5),
    .sum(pp_2_42_6),
    .cout(pp_2_43_1)
  );

  MG_FA fa_1_42_2(
    .a(pp_1_42_6),
    .b(pp_1_42_7),
    .cin(pp_1_42_8),
    .sum(pp_2_42_7),
    .cout(pp_2_43_2)
  );

  MG_FA fa_1_42_3(
    .a(pp_1_42_9),
    .b(pp_1_42_10),
    .cin(pp_1_42_11),
    .sum(pp_2_42_8),
    .cout(pp_2_43_3)
  );

  assign pp_2_42_9 = pp_1_42_12;
  MG_FA fa_1_43_0(
    .a(pp_1_43_0),
    .b(pp_1_43_1),
    .cin(pp_1_43_2),
    .sum(pp_2_43_4),
    .cout(pp_2_44_0)
  );

  MG_FA fa_1_43_1(
    .a(pp_1_43_3),
    .b(pp_1_43_4),
    .cin(pp_1_43_5),
    .sum(pp_2_43_5),
    .cout(pp_2_44_1)
  );

  MG_FA fa_1_43_2(
    .a(pp_1_43_6),
    .b(pp_1_43_7),
    .cin(pp_1_43_8),
    .sum(pp_2_43_6),
    .cout(pp_2_44_2)
  );

  MG_FA fa_1_43_3(
    .a(pp_1_43_9),
    .b(pp_1_43_10),
    .cin(pp_1_43_11),
    .sum(pp_2_43_7),
    .cout(pp_2_44_3)
  );

  MG_FA fa_1_43_4(
    .a(pp_1_43_12),
    .b(pp_1_43_13),
    .cin(pp_1_43_14),
    .sum(pp_2_43_8),
    .cout(pp_2_44_4)
  );

  MG_FA fa_1_44_0(
    .a(pp_1_44_0),
    .b(pp_1_44_1),
    .cin(pp_1_44_2),
    .sum(pp_2_44_5),
    .cout(pp_2_45_0)
  );

  MG_FA fa_1_44_1(
    .a(pp_1_44_3),
    .b(pp_1_44_4),
    .cin(pp_1_44_5),
    .sum(pp_2_44_6),
    .cout(pp_2_45_1)
  );

  MG_FA fa_1_44_2(
    .a(pp_1_44_6),
    .b(pp_1_44_7),
    .cin(pp_1_44_8),
    .sum(pp_2_44_7),
    .cout(pp_2_45_2)
  );

  MG_FA fa_1_44_3(
    .a(pp_1_44_9),
    .b(pp_1_44_10),
    .cin(pp_1_44_11),
    .sum(pp_2_44_8),
    .cout(pp_2_45_3)
  );

  MG_FA fa_1_44_4(
    .a(pp_1_44_12),
    .b(pp_1_44_13),
    .cin(pp_1_44_14),
    .sum(pp_2_44_9),
    .cout(pp_2_45_4)
  );

  MG_FA fa_1_44_5(
    .a(pp_1_44_15),
    .b(pp_1_44_16),
    .cin(pp_1_44_17),
    .sum(pp_2_44_10),
    .cout(pp_2_45_5)
  );

  MG_FA fa_1_44_6(
    .a(pp_1_44_18),
    .b(pp_1_44_19),
    .cin(pp_1_44_20),
    .sum(pp_2_44_11),
    .cout(pp_2_45_6)
  );

  assign pp_2_44_12 = pp_1_44_21;
  assign pp_2_44_13 = pp_1_44_22;
  assign pp_2_44_14 = pp_1_44_23;
  assign pp_2_44_15 = pp_1_44_24;
  MG_FA fa_1_45_0(
    .a(pp_1_45_0),
    .b(pp_1_45_1),
    .cin(pp_1_45_2),
    .sum(pp_2_45_7),
    .cout(pp_2_46_0)
  );

  MG_FA fa_1_45_1(
    .a(pp_1_45_3),
    .b(pp_1_45_4),
    .cin(pp_1_45_5),
    .sum(pp_2_45_8),
    .cout(pp_2_46_1)
  );

  MG_FA fa_1_46_0(
    .a(pp_1_46_0),
    .b(pp_1_46_1),
    .cin(pp_1_46_2),
    .sum(pp_2_46_2),
    .cout(pp_2_47_0)
  );

  MG_FA fa_1_46_1(
    .a(pp_1_46_3),
    .b(pp_1_46_4),
    .cin(pp_1_46_5),
    .sum(pp_2_46_3),
    .cout(pp_2_47_1)
  );

  MG_FA fa_1_46_2(
    .a(pp_1_46_6),
    .b(pp_1_46_7),
    .cin(pp_1_46_8),
    .sum(pp_2_46_4),
    .cout(pp_2_47_2)
  );

  MG_FA fa_1_46_3(
    .a(pp_1_46_9),
    .b(pp_1_46_10),
    .cin(pp_1_46_11),
    .sum(pp_2_46_5),
    .cout(pp_2_47_3)
  );

  MG_FA fa_1_46_4(
    .a(pp_1_46_12),
    .b(pp_1_46_13),
    .cin(pp_1_46_14),
    .sum(pp_2_46_6),
    .cout(pp_2_47_4)
  );

  MG_FA fa_1_47_0(
    .a(pp_1_47_0),
    .b(pp_1_47_1),
    .cin(pp_1_47_2),
    .sum(pp_2_47_5),
    .cout(pp_2_48_0)
  );

  MG_FA fa_1_47_1(
    .a(pp_1_47_3),
    .b(pp_1_47_4),
    .cin(pp_1_47_5),
    .sum(pp_2_47_6),
    .cout(pp_2_48_1)
  );

  MG_FA fa_1_47_2(
    .a(pp_1_47_6),
    .b(pp_1_47_7),
    .cin(pp_1_47_8),
    .sum(pp_2_47_7),
    .cout(pp_2_48_2)
  );

  MG_FA fa_1_47_3(
    .a(pp_1_47_9),
    .b(pp_1_47_10),
    .cin(pp_1_47_11),
    .sum(pp_2_47_8),
    .cout(pp_2_48_3)
  );

  MG_FA fa_1_48_0(
    .a(pp_1_48_0),
    .b(pp_1_48_1),
    .cin(pp_1_48_2),
    .sum(pp_2_48_4),
    .cout(pp_2_49_0)
  );

  MG_FA fa_1_48_1(
    .a(pp_1_48_3),
    .b(pp_1_48_4),
    .cin(pp_1_48_5),
    .sum(pp_2_48_5),
    .cout(pp_2_49_1)
  );

  MG_FA fa_1_48_2(
    .a(pp_1_48_6),
    .b(pp_1_48_7),
    .cin(pp_1_48_8),
    .sum(pp_2_48_6),
    .cout(pp_2_49_2)
  );

  MG_FA fa_1_49_0(
    .a(pp_1_49_0),
    .b(pp_1_49_1),
    .cin(pp_1_49_2),
    .sum(pp_2_49_3),
    .cout(pp_2_50_0)
  );

  MG_FA fa_1_49_1(
    .a(pp_1_49_3),
    .b(pp_1_49_4),
    .cin(pp_1_49_5),
    .sum(pp_2_49_4),
    .cout(pp_2_50_1)
  );

  MG_FA fa_1_49_2(
    .a(pp_1_49_6),
    .b(pp_1_49_7),
    .cin(pp_1_49_8),
    .sum(pp_2_49_5),
    .cout(pp_2_50_2)
  );

  assign pp_2_49_6 = pp_1_49_9;
  assign pp_2_49_7 = pp_1_49_10;
  MG_FA fa_1_50_0(
    .a(pp_1_50_0),
    .b(pp_1_50_1),
    .cin(pp_1_50_2),
    .sum(pp_2_50_3),
    .cout(pp_2_51_0)
  );

  MG_FA fa_1_50_1(
    .a(pp_1_50_3),
    .b(pp_1_50_4),
    .cin(pp_1_50_5),
    .sum(pp_2_50_4),
    .cout(pp_2_51_1)
  );

  MG_FA fa_1_50_2(
    .a(pp_1_50_6),
    .b(pp_1_50_7),
    .cin(pp_1_50_8),
    .sum(pp_2_50_5),
    .cout(pp_2_51_2)
  );

  MG_FA fa_1_51_0(
    .a(pp_1_51_0),
    .b(pp_1_51_1),
    .cin(pp_1_51_2),
    .sum(pp_2_51_3),
    .cout(pp_2_52_0)
  );

  MG_FA fa_1_51_1(
    .a(pp_1_51_3),
    .b(pp_1_51_4),
    .cin(pp_1_51_5),
    .sum(pp_2_51_4),
    .cout(pp_2_52_1)
  );

  assign pp_2_51_5 = pp_1_51_6;
  assign pp_2_51_6 = pp_1_51_7;
  MG_FA fa_1_52_0(
    .a(pp_1_52_0),
    .b(pp_1_52_1),
    .cin(pp_1_52_2),
    .sum(pp_2_52_2),
    .cout(pp_2_53_0)
  );

  MG_FA fa_1_52_1(
    .a(pp_1_52_3),
    .b(pp_1_52_4),
    .cin(pp_1_52_5),
    .sum(pp_2_52_3),
    .cout(pp_2_53_1)
  );

  MG_FA fa_1_52_2(
    .a(pp_1_52_6),
    .b(pp_1_52_7),
    .cin(pp_1_52_8),
    .sum(pp_2_52_4),
    .cout(pp_2_53_2)
  );

  MG_FA fa_1_53_0(
    .a(pp_1_53_0),
    .b(pp_1_53_1),
    .cin(pp_1_53_2),
    .sum(pp_2_53_3),
    .cout(pp_2_54_0)
  );

  MG_FA fa_1_53_1(
    .a(pp_1_53_3),
    .b(pp_1_53_4),
    .cin(pp_1_53_5),
    .sum(pp_2_53_4),
    .cout(pp_2_54_1)
  );

  assign pp_2_53_5 = pp_1_53_6;
  MG_FA fa_1_54_0(
    .a(pp_1_54_0),
    .b(pp_1_54_1),
    .cin(pp_1_54_2),
    .sum(pp_2_54_2),
    .cout(pp_2_55_0)
  );

  MG_FA fa_1_54_1(
    .a(pp_1_54_3),
    .b(pp_1_54_4),
    .cin(pp_1_54_5),
    .sum(pp_2_54_3),
    .cout(pp_2_55_1)
  );

  MG_FA fa_1_55_0(
    .a(pp_1_55_0),
    .b(pp_1_55_1),
    .cin(pp_1_55_2),
    .sum(pp_2_55_2),
    .cout(pp_2_56_0)
  );

  MG_FA fa_1_55_1(
    .a(pp_1_55_3),
    .b(pp_1_55_4),
    .cin(pp_1_55_5),
    .sum(pp_2_55_3),
    .cout(pp_2_56_1)
  );

  assign pp_2_55_4 = pp_1_55_6;
  MG_FA fa_1_56_0(
    .a(pp_1_56_0),
    .b(pp_1_56_1),
    .cin(pp_1_56_2),
    .sum(pp_2_56_2),
    .cout(pp_2_57_0)
  );

  MG_FA fa_1_56_1(
    .a(pp_1_56_3),
    .b(pp_1_56_4),
    .cin(pp_1_56_5),
    .sum(pp_2_56_3),
    .cout(pp_2_57_1)
  );

  MG_FA fa_1_56_2(
    .a(pp_1_56_6),
    .b(pp_1_56_7),
    .cin(pp_1_56_8),
    .sum(pp_2_56_4),
    .cout(pp_2_57_2)
  );

  assign pp_2_57_3 = pp_1_57_0;
  assign pp_2_57_4 = pp_1_57_1;
  MG_FA fa_1_58_0(
    .a(pp_1_58_0),
    .b(pp_1_58_1),
    .cin(pp_1_58_2),
    .sum(pp_2_58_0),
    .cout(pp_2_59_0)
  );

  MG_FA fa_1_58_1(
    .a(pp_1_58_3),
    .b(pp_1_58_4),
    .cin(pp_1_58_5),
    .sum(pp_2_58_1),
    .cout(pp_2_59_1)
  );

  assign pp_2_58_2 = pp_1_58_6;
  assign pp_2_59_2 = pp_1_59_0;
  assign pp_2_59_3 = pp_1_59_1;
  assign pp_2_59_4 = pp_1_59_2;
  assign pp_2_59_5 = pp_1_59_3;
  assign pp_2_60_0 = pp_1_60_0;
  assign pp_2_61_0 = pp_1_61_0;
  assign pp_2_61_1 = pp_1_61_1;
  assign pp_2_61_2 = pp_1_61_2;
  assign pp_2_62_0 = pp_1_62_0;
  assign pp_3_0_0 = pp_2_0_0;
  assign pp_3_1_0 = pp_2_1_0;
  assign pp_3_1_1 = pp_2_1_1;
  assign pp_3_2_0 = pp_2_2_0;
  assign pp_3_2_1 = pp_2_2_1;
  assign pp_3_2_2 = pp_2_2_2;
  MG_HA ha_2_3_0(
    .a(pp_2_3_0),
    .b(pp_2_3_1),
    .sum(pp_3_3_0),
    .cout(pp_3_4_0)
  );

  assign pp_3_3_1 = pp_2_3_2;
  assign pp_3_3_2 = pp_2_3_3;
  MG_FA fa_2_4_0(
    .a(pp_2_4_0),
    .b(pp_2_4_1),
    .cin(pp_2_4_2),
    .sum(pp_3_4_1),
    .cout(pp_3_5_0)
  );

  MG_FA fa_2_5_0(
    .a(pp_2_5_0),
    .b(pp_2_5_1),
    .cin(pp_2_5_2),
    .sum(pp_3_5_1),
    .cout(pp_3_6_0)
  );

  MG_FA fa_2_6_0(
    .a(pp_2_6_0),
    .b(pp_2_6_1),
    .cin(pp_2_6_2),
    .sum(pp_3_6_1),
    .cout(pp_3_7_0)
  );

  MG_FA fa_2_6_1(
    .a(pp_2_6_3),
    .b(pp_2_6_4),
    .cin(pp_2_6_5),
    .sum(pp_3_6_2),
    .cout(pp_3_7_1)
  );

  assign pp_3_6_3 = pp_2_6_6;
  assign pp_3_7_2 = pp_2_7_0;
  assign pp_3_7_3 = pp_2_7_1;
  assign pp_3_8_0 = pp_2_8_0;
  assign pp_3_8_1 = pp_2_8_1;
  assign pp_3_8_2 = pp_2_8_2;
  assign pp_3_8_3 = pp_2_8_3;
  assign pp_3_8_4 = pp_2_8_4;
  assign pp_3_8_5 = pp_2_8_5;
  MG_FA fa_2_9_0(
    .a(pp_2_9_0),
    .b(pp_2_9_1),
    .cin(pp_2_9_2),
    .sum(pp_3_9_0),
    .cout(pp_3_10_0)
  );

  MG_FA fa_2_9_1(
    .a(pp_2_9_3),
    .b(pp_2_9_4),
    .cin(pp_2_9_5),
    .sum(pp_3_9_1),
    .cout(pp_3_10_1)
  );

  MG_FA fa_2_9_2(
    .a(pp_2_9_6),
    .b(pp_2_9_7),
    .cin(pp_2_9_8),
    .sum(pp_3_9_2),
    .cout(pp_3_10_2)
  );

  MG_FA fa_2_10_0(
    .a(pp_2_10_0),
    .b(pp_2_10_1),
    .cin(pp_2_10_2),
    .sum(pp_3_10_3),
    .cout(pp_3_11_0)
  );

  assign pp_3_10_4 = pp_2_10_3;
  MG_FA fa_2_11_0(
    .a(pp_2_11_0),
    .b(pp_2_11_1),
    .cin(pp_2_11_2),
    .sum(pp_3_11_1),
    .cout(pp_3_12_0)
  );

  MG_FA fa_2_11_1(
    .a(pp_2_11_3),
    .b(pp_2_11_4),
    .cin(pp_2_11_5),
    .sum(pp_3_11_2),
    .cout(pp_3_12_1)
  );

  assign pp_3_11_3 = pp_2_11_6;
  assign pp_3_11_4 = pp_2_11_7;
  assign pp_3_11_5 = pp_2_11_8;
  MG_FA fa_2_12_0(
    .a(pp_2_12_0),
    .b(pp_2_12_1),
    .cin(pp_2_12_2),
    .sum(pp_3_12_2),
    .cout(pp_3_13_0)
  );

  MG_FA fa_2_13_0(
    .a(pp_2_13_0),
    .b(pp_2_13_1),
    .cin(pp_2_13_2),
    .sum(pp_3_13_1),
    .cout(pp_3_14_0)
  );

  MG_FA fa_2_13_1(
    .a(pp_2_13_3),
    .b(pp_2_13_4),
    .cin(pp_2_13_5),
    .sum(pp_3_13_2),
    .cout(pp_3_14_1)
  );

  MG_FA fa_2_14_0(
    .a(pp_2_14_0),
    .b(pp_2_14_1),
    .cin(pp_2_14_2),
    .sum(pp_3_14_2),
    .cout(pp_3_15_0)
  );

  MG_FA fa_2_14_1(
    .a(pp_2_14_3),
    .b(pp_2_14_4),
    .cin(pp_2_14_5),
    .sum(pp_3_14_3),
    .cout(pp_3_15_1)
  );

  MG_FA fa_2_14_2(
    .a(pp_2_14_6),
    .b(pp_2_14_7),
    .cin(pp_2_14_8),
    .sum(pp_3_14_4),
    .cout(pp_3_15_2)
  );

  assign pp_3_14_5 = pp_2_14_9;
  assign pp_3_14_6 = pp_2_14_10;
  assign pp_3_14_7 = pp_2_14_11;
  assign pp_3_14_8 = pp_2_14_12;
  MG_FA fa_2_15_0(
    .a(pp_2_15_0),
    .b(pp_2_15_1),
    .cin(pp_2_15_2),
    .sum(pp_3_15_3),
    .cout(pp_3_16_0)
  );

  assign pp_3_15_4 = pp_2_15_3;
  assign pp_3_16_1 = pp_2_16_0;
  assign pp_3_16_2 = pp_2_16_1;
  assign pp_3_16_3 = pp_2_16_2;
  assign pp_3_16_4 = pp_2_16_3;
  assign pp_3_16_5 = pp_2_16_4;
  assign pp_3_16_6 = pp_2_16_5;
  assign pp_3_16_7 = pp_2_16_6;
  assign pp_3_16_8 = pp_2_16_7;
  MG_FA fa_2_17_0(
    .a(pp_2_17_0),
    .b(pp_2_17_1),
    .cin(pp_2_17_2),
    .sum(pp_3_17_0),
    .cout(pp_3_18_0)
  );

  MG_FA fa_2_17_1(
    .a(pp_2_17_3),
    .b(pp_2_17_4),
    .cin(pp_2_17_5),
    .sum(pp_3_17_1),
    .cout(pp_3_18_1)
  );

  MG_FA fa_2_17_2(
    .a(pp_2_17_6),
    .b(pp_2_17_7),
    .cin(pp_2_17_8),
    .sum(pp_3_17_2),
    .cout(pp_3_18_2)
  );

  assign pp_3_18_3 = pp_2_18_0;
  assign pp_3_18_4 = pp_2_18_1;
  assign pp_3_18_5 = pp_2_18_2;
  assign pp_3_18_6 = pp_2_18_3;
  assign pp_3_18_7 = pp_2_18_4;
  assign pp_3_18_8 = pp_2_18_5;
  assign pp_3_18_9 = pp_2_18_6;
  assign pp_3_18_10 = pp_2_18_7;
  MG_FA fa_2_19_0(
    .a(pp_2_19_0),
    .b(pp_2_19_1),
    .cin(pp_2_19_2),
    .sum(pp_3_19_0),
    .cout(pp_3_20_0)
  );

  MG_FA fa_2_19_1(
    .a(pp_2_19_3),
    .b(pp_2_19_4),
    .cin(pp_2_19_5),
    .sum(pp_3_19_1),
    .cout(pp_3_20_1)
  );

  MG_FA fa_2_19_2(
    .a(pp_2_19_6),
    .b(pp_2_19_7),
    .cin(pp_2_19_8),
    .sum(pp_3_19_2),
    .cout(pp_3_20_2)
  );

  MG_FA fa_2_20_0(
    .a(pp_2_20_0),
    .b(pp_2_20_1),
    .cin(pp_2_20_2),
    .sum(pp_3_20_3),
    .cout(pp_3_21_0)
  );

  MG_FA fa_2_20_1(
    .a(pp_2_20_3),
    .b(pp_2_20_4),
    .cin(pp_2_20_5),
    .sum(pp_3_20_4),
    .cout(pp_3_21_1)
  );

  MG_FA fa_2_20_2(
    .a(pp_2_20_6),
    .b(pp_2_20_7),
    .cin(pp_2_20_8),
    .sum(pp_3_20_5),
    .cout(pp_3_21_2)
  );

  MG_FA fa_2_21_0(
    .a(pp_2_21_0),
    .b(pp_2_21_1),
    .cin(pp_2_21_2),
    .sum(pp_3_21_3),
    .cout(pp_3_22_0)
  );

  MG_FA fa_2_21_1(
    .a(pp_2_21_3),
    .b(pp_2_21_4),
    .cin(pp_2_21_5),
    .sum(pp_3_21_4),
    .cout(pp_3_22_1)
  );

  assign pp_3_21_5 = pp_2_21_6;
  assign pp_3_21_6 = pp_2_21_7;
  assign pp_3_21_7 = pp_2_21_8;
  assign pp_3_21_8 = pp_2_21_9;
  MG_FA fa_2_22_0(
    .a(pp_2_22_0),
    .b(pp_2_22_1),
    .cin(pp_2_22_2),
    .sum(pp_3_22_2),
    .cout(pp_3_23_0)
  );

  MG_FA fa_2_22_1(
    .a(pp_2_22_3),
    .b(pp_2_22_4),
    .cin(pp_2_22_5),
    .sum(pp_3_22_3),
    .cout(pp_3_23_1)
  );

  MG_FA fa_2_22_2(
    .a(pp_2_22_6),
    .b(pp_2_22_7),
    .cin(pp_2_22_8),
    .sum(pp_3_22_4),
    .cout(pp_3_23_2)
  );

  MG_FA fa_2_22_3(
    .a(pp_2_22_9),
    .b(pp_2_22_10),
    .cin(pp_2_22_11),
    .sum(pp_3_22_5),
    .cout(pp_3_23_3)
  );

  MG_FA fa_2_22_4(
    .a(pp_2_22_12),
    .b(pp_2_22_13),
    .cin(pp_2_22_14),
    .sum(pp_3_22_6),
    .cout(pp_3_23_4)
  );

  MG_FA fa_2_22_5(
    .a(pp_2_22_15),
    .b(pp_2_22_16),
    .cin(pp_2_22_17),
    .sum(pp_3_22_7),
    .cout(pp_3_23_5)
  );

  assign pp_3_22_8 = pp_2_22_18;
  assign pp_3_22_9 = pp_2_22_19;
  assign pp_3_22_10 = pp_2_22_20;
  MG_FA fa_2_23_0(
    .a(pp_2_23_0),
    .b(pp_2_23_1),
    .cin(pp_2_23_2),
    .sum(pp_3_23_6),
    .cout(pp_3_24_0)
  );

  assign pp_3_23_7 = pp_2_23_3;
  assign pp_3_23_8 = pp_2_23_4;
  MG_FA fa_2_24_0(
    .a(pp_2_24_0),
    .b(pp_2_24_1),
    .cin(pp_2_24_2),
    .sum(pp_3_24_1),
    .cout(pp_3_25_0)
  );

  MG_FA fa_2_24_1(
    .a(pp_2_24_3),
    .b(pp_2_24_4),
    .cin(pp_2_24_5),
    .sum(pp_3_24_2),
    .cout(pp_3_25_1)
  );

  MG_FA fa_2_24_2(
    .a(pp_2_24_6),
    .b(pp_2_24_7),
    .cin(pp_2_24_8),
    .sum(pp_3_24_3),
    .cout(pp_3_25_2)
  );

  MG_FA fa_2_24_3(
    .a(pp_2_24_9),
    .b(pp_2_24_10),
    .cin(pp_2_24_11),
    .sum(pp_3_24_4),
    .cout(pp_3_25_3)
  );

  MG_FA fa_2_25_0(
    .a(pp_2_25_0),
    .b(pp_2_25_1),
    .cin(pp_2_25_2),
    .sum(pp_3_25_4),
    .cout(pp_3_26_0)
  );

  MG_FA fa_2_25_1(
    .a(pp_2_25_3),
    .b(pp_2_25_4),
    .cin(pp_2_25_5),
    .sum(pp_3_25_5),
    .cout(pp_3_26_1)
  );

  MG_FA fa_2_25_2(
    .a(pp_2_25_6),
    .b(pp_2_25_7),
    .cin(pp_2_25_8),
    .sum(pp_3_25_6),
    .cout(pp_3_26_2)
  );

  assign pp_3_25_7 = pp_2_25_9;
  assign pp_3_25_8 = pp_2_25_10;
  assign pp_3_25_9 = pp_2_25_11;
  assign pp_3_25_10 = pp_2_25_12;
  assign pp_3_25_11 = pp_2_25_13;
  assign pp_3_25_12 = pp_2_25_14;
  assign pp_3_25_13 = pp_2_25_15;
  assign pp_3_25_14 = pp_2_25_16;
  MG_FA fa_2_26_0(
    .a(pp_2_26_0),
    .b(pp_2_26_1),
    .cin(pp_2_26_2),
    .sum(pp_3_26_3),
    .cout(pp_3_27_0)
  );

  MG_FA fa_2_26_1(
    .a(pp_2_26_3),
    .b(pp_2_26_4),
    .cin(pp_2_26_5),
    .sum(pp_3_26_4),
    .cout(pp_3_27_1)
  );

  MG_FA fa_2_26_2(
    .a(pp_2_26_6),
    .b(pp_2_26_7),
    .cin(pp_2_26_8),
    .sum(pp_3_26_5),
    .cout(pp_3_27_2)
  );

  MG_FA fa_2_26_3(
    .a(pp_2_26_9),
    .b(pp_2_26_10),
    .cin(pp_2_26_11),
    .sum(pp_3_26_6),
    .cout(pp_3_27_3)
  );

  MG_FA fa_2_26_4(
    .a(pp_2_26_12),
    .b(pp_2_26_13),
    .cin(pp_2_26_14),
    .sum(pp_3_26_7),
    .cout(pp_3_27_4)
  );

  MG_FA fa_2_27_0(
    .a(pp_2_27_0),
    .b(pp_2_27_1),
    .cin(pp_2_27_2),
    .sum(pp_3_27_5),
    .cout(pp_3_28_0)
  );

  MG_FA fa_2_27_1(
    .a(pp_2_27_3),
    .b(pp_2_27_4),
    .cin(pp_2_27_5),
    .sum(pp_3_27_6),
    .cout(pp_3_28_1)
  );

  MG_FA fa_2_27_2(
    .a(pp_2_27_6),
    .b(pp_2_27_7),
    .cin(pp_2_27_8),
    .sum(pp_3_27_7),
    .cout(pp_3_28_2)
  );

  MG_FA fa_2_27_3(
    .a(pp_2_27_9),
    .b(pp_2_27_10),
    .cin(pp_2_27_11),
    .sum(pp_3_27_8),
    .cout(pp_3_28_3)
  );

  MG_FA fa_2_28_0(
    .a(pp_2_28_0),
    .b(pp_2_28_1),
    .cin(pp_2_28_2),
    .sum(pp_3_28_4),
    .cout(pp_3_29_0)
  );

  MG_FA fa_2_28_1(
    .a(pp_2_28_3),
    .b(pp_2_28_4),
    .cin(pp_2_28_5),
    .sum(pp_3_28_5),
    .cout(pp_3_29_1)
  );

  MG_FA fa_2_28_2(
    .a(pp_2_28_6),
    .b(pp_2_28_7),
    .cin(pp_2_28_8),
    .sum(pp_3_28_6),
    .cout(pp_3_29_2)
  );

  MG_FA fa_2_28_3(
    .a(pp_2_28_9),
    .b(pp_2_28_10),
    .cin(pp_2_28_11),
    .sum(pp_3_28_7),
    .cout(pp_3_29_3)
  );

  assign pp_3_28_8 = pp_2_28_12;
  MG_FA fa_2_29_0(
    .a(pp_2_29_0),
    .b(pp_2_29_1),
    .cin(pp_2_29_2),
    .sum(pp_3_29_4),
    .cout(pp_3_30_0)
  );

  MG_FA fa_2_29_1(
    .a(pp_2_29_3),
    .b(pp_2_29_4),
    .cin(pp_2_29_5),
    .sum(pp_3_29_5),
    .cout(pp_3_30_1)
  );

  MG_FA fa_2_29_2(
    .a(pp_2_29_6),
    .b(pp_2_29_7),
    .cin(pp_2_29_8),
    .sum(pp_3_29_6),
    .cout(pp_3_30_2)
  );

  MG_FA fa_2_29_3(
    .a(pp_2_29_9),
    .b(pp_2_29_10),
    .cin(pp_2_29_11),
    .sum(pp_3_29_7),
    .cout(pp_3_30_3)
  );

  assign pp_3_29_8 = pp_2_29_12;
  MG_FA fa_2_30_0(
    .a(pp_2_30_0),
    .b(pp_2_30_1),
    .cin(pp_2_30_2),
    .sum(pp_3_30_4),
    .cout(pp_3_31_0)
  );

  MG_FA fa_2_30_1(
    .a(pp_2_30_3),
    .b(pp_2_30_4),
    .cin(pp_2_30_5),
    .sum(pp_3_30_5),
    .cout(pp_3_31_1)
  );

  MG_FA fa_2_30_2(
    .a(pp_2_30_6),
    .b(pp_2_30_7),
    .cin(pp_2_30_8),
    .sum(pp_3_30_6),
    .cout(pp_3_31_2)
  );

  MG_FA fa_2_30_3(
    .a(pp_2_30_9),
    .b(pp_2_30_10),
    .cin(pp_2_30_11),
    .sum(pp_3_30_7),
    .cout(pp_3_31_3)
  );

  assign pp_3_30_8 = pp_2_30_12;
  MG_FA fa_2_31_0(
    .a(pp_2_31_0),
    .b(pp_2_31_1),
    .cin(pp_2_31_2),
    .sum(pp_3_31_4),
    .cout(pp_3_32_0)
  );

  MG_FA fa_2_31_1(
    .a(pp_2_31_3),
    .b(pp_2_31_4),
    .cin(pp_2_31_5),
    .sum(pp_3_31_5),
    .cout(pp_3_32_1)
  );

  MG_FA fa_2_31_2(
    .a(pp_2_31_6),
    .b(pp_2_31_7),
    .cin(pp_2_31_8),
    .sum(pp_3_31_6),
    .cout(pp_3_32_2)
  );

  MG_FA fa_2_31_3(
    .a(pp_2_31_9),
    .b(pp_2_31_10),
    .cin(pp_2_31_11),
    .sum(pp_3_31_7),
    .cout(pp_3_32_3)
  );

  MG_FA fa_2_31_4(
    .a(pp_2_31_12),
    .b(pp_2_31_13),
    .cin(pp_2_31_14),
    .sum(pp_3_31_8),
    .cout(pp_3_32_4)
  );

  MG_FA fa_2_32_0(
    .a(pp_2_32_0),
    .b(pp_2_32_1),
    .cin(pp_2_32_2),
    .sum(pp_3_32_5),
    .cout(pp_3_33_0)
  );

  MG_FA fa_2_32_1(
    .a(pp_2_32_3),
    .b(pp_2_32_4),
    .cin(pp_2_32_5),
    .sum(pp_3_32_6),
    .cout(pp_3_33_1)
  );

  MG_FA fa_2_32_2(
    .a(pp_2_32_6),
    .b(pp_2_32_7),
    .cin(pp_2_32_8),
    .sum(pp_3_32_7),
    .cout(pp_3_33_2)
  );

  MG_FA fa_2_32_3(
    .a(pp_2_32_9),
    .b(pp_2_32_10),
    .cin(pp_2_32_11),
    .sum(pp_3_32_8),
    .cout(pp_3_33_3)
  );

  assign pp_3_32_9 = pp_2_32_12;
  assign pp_3_32_10 = pp_2_32_13;
  MG_FA fa_2_33_0(
    .a(pp_2_33_0),
    .b(pp_2_33_1),
    .cin(pp_2_33_2),
    .sum(pp_3_33_4),
    .cout(pp_3_34_0)
  );

  MG_FA fa_2_33_1(
    .a(pp_2_33_3),
    .b(pp_2_33_4),
    .cin(pp_2_33_5),
    .sum(pp_3_33_5),
    .cout(pp_3_34_1)
  );

  MG_FA fa_2_33_2(
    .a(pp_2_33_6),
    .b(pp_2_33_7),
    .cin(pp_2_33_8),
    .sum(pp_3_33_6),
    .cout(pp_3_34_2)
  );

  MG_FA fa_2_33_3(
    .a(pp_2_33_9),
    .b(pp_2_33_10),
    .cin(pp_2_33_11),
    .sum(pp_3_33_7),
    .cout(pp_3_34_3)
  );

  MG_FA fa_2_33_4(
    .a(pp_2_33_12),
    .b(pp_2_33_13),
    .cin(pp_2_33_14),
    .sum(pp_3_33_8),
    .cout(pp_3_34_4)
  );

  MG_FA fa_2_34_0(
    .a(pp_2_34_0),
    .b(pp_2_34_1),
    .cin(pp_2_34_2),
    .sum(pp_3_34_5),
    .cout(pp_3_35_0)
  );

  MG_FA fa_2_34_1(
    .a(pp_2_34_3),
    .b(pp_2_34_4),
    .cin(pp_2_34_5),
    .sum(pp_3_34_6),
    .cout(pp_3_35_1)
  );

  MG_FA fa_2_34_2(
    .a(pp_2_34_6),
    .b(pp_2_34_7),
    .cin(pp_2_34_8),
    .sum(pp_3_34_7),
    .cout(pp_3_35_2)
  );

  MG_FA fa_2_34_3(
    .a(pp_2_34_9),
    .b(pp_2_34_10),
    .cin(pp_2_34_11),
    .sum(pp_3_34_8),
    .cout(pp_3_35_3)
  );

  assign pp_3_34_9 = pp_2_34_12;
  MG_FA fa_2_35_0(
    .a(pp_2_35_0),
    .b(pp_2_35_1),
    .cin(pp_2_35_2),
    .sum(pp_3_35_4),
    .cout(pp_3_36_0)
  );

  MG_FA fa_2_35_1(
    .a(pp_2_35_3),
    .b(pp_2_35_4),
    .cin(pp_2_35_5),
    .sum(pp_3_35_5),
    .cout(pp_3_36_1)
  );

  MG_FA fa_2_35_2(
    .a(pp_2_35_6),
    .b(pp_2_35_7),
    .cin(pp_2_35_8),
    .sum(pp_3_35_6),
    .cout(pp_3_36_2)
  );

  MG_FA fa_2_35_3(
    .a(pp_2_35_9),
    .b(pp_2_35_10),
    .cin(pp_2_35_11),
    .sum(pp_3_35_7),
    .cout(pp_3_36_3)
  );

  assign pp_3_35_8 = pp_2_35_12;
  assign pp_3_35_9 = pp_2_35_13;
  MG_FA fa_2_36_0(
    .a(pp_2_36_0),
    .b(pp_2_36_1),
    .cin(pp_2_36_2),
    .sum(pp_3_36_4),
    .cout(pp_3_37_0)
  );

  MG_FA fa_2_36_1(
    .a(pp_2_36_3),
    .b(pp_2_36_4),
    .cin(pp_2_36_5),
    .sum(pp_3_36_5),
    .cout(pp_3_37_1)
  );

  MG_FA fa_2_36_2(
    .a(pp_2_36_6),
    .b(pp_2_36_7),
    .cin(pp_2_36_8),
    .sum(pp_3_36_6),
    .cout(pp_3_37_2)
  );

  MG_FA fa_2_36_3(
    .a(pp_2_36_9),
    .b(pp_2_36_10),
    .cin(pp_2_36_11),
    .sum(pp_3_36_7),
    .cout(pp_3_37_3)
  );

  MG_FA fa_2_37_0(
    .a(pp_2_37_0),
    .b(pp_2_37_1),
    .cin(pp_2_37_2),
    .sum(pp_3_37_4),
    .cout(pp_3_38_0)
  );

  MG_FA fa_2_37_1(
    .a(pp_2_37_3),
    .b(pp_2_37_4),
    .cin(pp_2_37_5),
    .sum(pp_3_37_5),
    .cout(pp_3_38_1)
  );

  MG_FA fa_2_37_2(
    .a(pp_2_37_6),
    .b(pp_2_37_7),
    .cin(pp_2_37_8),
    .sum(pp_3_37_6),
    .cout(pp_3_38_2)
  );

  MG_FA fa_2_37_3(
    .a(pp_2_37_9),
    .b(pp_2_37_10),
    .cin(pp_2_37_11),
    .sum(pp_3_37_7),
    .cout(pp_3_38_3)
  );

  assign pp_3_37_8 = pp_2_37_12;
  MG_FA fa_2_38_0(
    .a(pp_2_38_0),
    .b(pp_2_38_1),
    .cin(pp_2_38_2),
    .sum(pp_3_38_4),
    .cout(pp_3_39_0)
  );

  MG_FA fa_2_38_1(
    .a(pp_2_38_3),
    .b(pp_2_38_4),
    .cin(pp_2_38_5),
    .sum(pp_3_38_5),
    .cout(pp_3_39_1)
  );

  MG_FA fa_2_38_2(
    .a(pp_2_38_6),
    .b(pp_2_38_7),
    .cin(pp_2_38_8),
    .sum(pp_3_38_6),
    .cout(pp_3_39_2)
  );

  MG_FA fa_2_38_3(
    .a(pp_2_38_9),
    .b(pp_2_38_10),
    .cin(pp_2_38_11),
    .sum(pp_3_38_7),
    .cout(pp_3_39_3)
  );

  assign pp_3_38_8 = pp_2_38_12;
  MG_FA fa_2_39_0(
    .a(pp_2_39_0),
    .b(pp_2_39_1),
    .cin(pp_2_39_2),
    .sum(pp_3_39_4),
    .cout(pp_3_40_0)
  );

  MG_FA fa_2_39_1(
    .a(pp_2_39_3),
    .b(pp_2_39_4),
    .cin(pp_2_39_5),
    .sum(pp_3_39_5),
    .cout(pp_3_40_1)
  );

  MG_FA fa_2_39_2(
    .a(pp_2_39_6),
    .b(pp_2_39_7),
    .cin(pp_2_39_8),
    .sum(pp_3_39_6),
    .cout(pp_3_40_2)
  );

  assign pp_3_39_7 = pp_2_39_9;
  assign pp_3_39_8 = pp_2_39_10;
  MG_FA fa_2_40_0(
    .a(pp_2_40_0),
    .b(pp_2_40_1),
    .cin(pp_2_40_2),
    .sum(pp_3_40_3),
    .cout(pp_3_41_0)
  );

  MG_FA fa_2_40_1(
    .a(pp_2_40_3),
    .b(pp_2_40_4),
    .cin(pp_2_40_5),
    .sum(pp_3_40_4),
    .cout(pp_3_41_1)
  );

  MG_FA fa_2_40_2(
    .a(pp_2_40_6),
    .b(pp_2_40_7),
    .cin(pp_2_40_8),
    .sum(pp_3_40_5),
    .cout(pp_3_41_2)
  );

  MG_FA fa_2_40_3(
    .a(pp_2_40_9),
    .b(pp_2_40_10),
    .cin(pp_2_40_11),
    .sum(pp_3_40_6),
    .cout(pp_3_41_3)
  );

  MG_FA fa_2_41_0(
    .a(pp_2_41_0),
    .b(pp_2_41_1),
    .cin(pp_2_41_2),
    .sum(pp_3_41_4),
    .cout(pp_3_42_0)
  );

  MG_FA fa_2_41_1(
    .a(pp_2_41_3),
    .b(pp_2_41_4),
    .cin(pp_2_41_5),
    .sum(pp_3_41_5),
    .cout(pp_3_42_1)
  );

  assign pp_3_41_6 = pp_2_41_6;
  assign pp_3_41_7 = pp_2_41_7;
  assign pp_3_41_8 = pp_2_41_8;
  assign pp_3_41_9 = pp_2_41_9;
  assign pp_3_41_10 = pp_2_41_10;
  assign pp_3_41_11 = pp_2_41_11;
  MG_FA fa_2_42_0(
    .a(pp_2_42_0),
    .b(pp_2_42_1),
    .cin(pp_2_42_2),
    .sum(pp_3_42_2),
    .cout(pp_3_43_0)
  );

  MG_FA fa_2_42_1(
    .a(pp_2_42_3),
    .b(pp_2_42_4),
    .cin(pp_2_42_5),
    .sum(pp_3_42_3),
    .cout(pp_3_43_1)
  );

  MG_FA fa_2_42_2(
    .a(pp_2_42_6),
    .b(pp_2_42_7),
    .cin(pp_2_42_8),
    .sum(pp_3_42_4),
    .cout(pp_3_43_2)
  );

  assign pp_3_42_5 = pp_2_42_9;
  MG_FA fa_2_43_0(
    .a(pp_2_43_0),
    .b(pp_2_43_1),
    .cin(pp_2_43_2),
    .sum(pp_3_43_3),
    .cout(pp_3_44_0)
  );

  MG_FA fa_2_43_1(
    .a(pp_2_43_3),
    .b(pp_2_43_4),
    .cin(pp_2_43_5),
    .sum(pp_3_43_4),
    .cout(pp_3_44_1)
  );

  MG_FA fa_2_43_2(
    .a(pp_2_43_6),
    .b(pp_2_43_7),
    .cin(pp_2_43_8),
    .sum(pp_3_43_5),
    .cout(pp_3_44_2)
  );

  MG_FA fa_2_44_0(
    .a(pp_2_44_0),
    .b(pp_2_44_1),
    .cin(pp_2_44_2),
    .sum(pp_3_44_3),
    .cout(pp_3_45_0)
  );

  MG_FA fa_2_44_1(
    .a(pp_2_44_3),
    .b(pp_2_44_4),
    .cin(pp_2_44_5),
    .sum(pp_3_44_4),
    .cout(pp_3_45_1)
  );

  MG_FA fa_2_44_2(
    .a(pp_2_44_6),
    .b(pp_2_44_7),
    .cin(pp_2_44_8),
    .sum(pp_3_44_5),
    .cout(pp_3_45_2)
  );

  MG_FA fa_2_44_3(
    .a(pp_2_44_9),
    .b(pp_2_44_10),
    .cin(pp_2_44_11),
    .sum(pp_3_44_6),
    .cout(pp_3_45_3)
  );

  MG_FA fa_2_44_4(
    .a(pp_2_44_12),
    .b(pp_2_44_13),
    .cin(pp_2_44_14),
    .sum(pp_3_44_7),
    .cout(pp_3_45_4)
  );

  assign pp_3_44_8 = pp_2_44_15;
  MG_FA fa_2_45_0(
    .a(pp_2_45_0),
    .b(pp_2_45_1),
    .cin(pp_2_45_2),
    .sum(pp_3_45_5),
    .cout(pp_3_46_0)
  );

  MG_FA fa_2_45_1(
    .a(pp_2_45_3),
    .b(pp_2_45_4),
    .cin(pp_2_45_5),
    .sum(pp_3_45_6),
    .cout(pp_3_46_1)
  );

  assign pp_3_45_7 = pp_2_45_6;
  assign pp_3_45_8 = pp_2_45_7;
  assign pp_3_45_9 = pp_2_45_8;
  assign pp_3_46_2 = pp_2_46_0;
  assign pp_3_46_3 = pp_2_46_1;
  assign pp_3_46_4 = pp_2_46_2;
  assign pp_3_46_5 = pp_2_46_3;
  assign pp_3_46_6 = pp_2_46_4;
  assign pp_3_46_7 = pp_2_46_5;
  assign pp_3_46_8 = pp_2_46_6;
  MG_FA fa_2_47_0(
    .a(pp_2_47_0),
    .b(pp_2_47_1),
    .cin(pp_2_47_2),
    .sum(pp_3_47_0),
    .cout(pp_3_48_0)
  );

  MG_FA fa_2_47_1(
    .a(pp_2_47_3),
    .b(pp_2_47_4),
    .cin(pp_2_47_5),
    .sum(pp_3_47_1),
    .cout(pp_3_48_1)
  );

  MG_FA fa_2_47_2(
    .a(pp_2_47_6),
    .b(pp_2_47_7),
    .cin(pp_2_47_8),
    .sum(pp_3_47_2),
    .cout(pp_3_48_2)
  );

  MG_FA fa_2_48_0(
    .a(pp_2_48_0),
    .b(pp_2_48_1),
    .cin(pp_2_48_2),
    .sum(pp_3_48_3),
    .cout(pp_3_49_0)
  );

  MG_FA fa_2_48_1(
    .a(pp_2_48_3),
    .b(pp_2_48_4),
    .cin(pp_2_48_5),
    .sum(pp_3_48_4),
    .cout(pp_3_49_1)
  );

  assign pp_3_48_5 = pp_2_48_6;
  MG_FA fa_2_49_0(
    .a(pp_2_49_0),
    .b(pp_2_49_1),
    .cin(pp_2_49_2),
    .sum(pp_3_49_2),
    .cout(pp_3_50_0)
  );

  MG_FA fa_2_49_1(
    .a(pp_2_49_3),
    .b(pp_2_49_4),
    .cin(pp_2_49_5),
    .sum(pp_3_49_3),
    .cout(pp_3_50_1)
  );

  assign pp_3_49_4 = pp_2_49_6;
  assign pp_3_49_5 = pp_2_49_7;
  MG_FA fa_2_50_0(
    .a(pp_2_50_0),
    .b(pp_2_50_1),
    .cin(pp_2_50_2),
    .sum(pp_3_50_2),
    .cout(pp_3_51_0)
  );

  assign pp_3_50_3 = pp_2_50_3;
  assign pp_3_50_4 = pp_2_50_4;
  assign pp_3_50_5 = pp_2_50_5;
  MG_FA fa_2_51_0(
    .a(pp_2_51_0),
    .b(pp_2_51_1),
    .cin(pp_2_51_2),
    .sum(pp_3_51_1),
    .cout(pp_3_52_0)
  );

  assign pp_3_51_2 = pp_2_51_3;
  assign pp_3_51_3 = pp_2_51_4;
  assign pp_3_51_4 = pp_2_51_5;
  assign pp_3_51_5 = pp_2_51_6;
  MG_FA fa_2_52_0(
    .a(pp_2_52_0),
    .b(pp_2_52_1),
    .cin(pp_2_52_2),
    .sum(pp_3_52_1),
    .cout(pp_3_53_0)
  );

  assign pp_3_52_2 = pp_2_52_3;
  assign pp_3_52_3 = pp_2_52_4;
  MG_FA fa_2_53_0(
    .a(pp_2_53_0),
    .b(pp_2_53_1),
    .cin(pp_2_53_2),
    .sum(pp_3_53_1),
    .cout(pp_3_54_0)
  );

  MG_FA fa_2_53_1(
    .a(pp_2_53_3),
    .b(pp_2_53_4),
    .cin(pp_2_53_5),
    .sum(pp_3_53_2),
    .cout(pp_3_54_1)
  );

  assign pp_3_54_2 = pp_2_54_0;
  assign pp_3_54_3 = pp_2_54_1;
  assign pp_3_54_4 = pp_2_54_2;
  assign pp_3_54_5 = pp_2_54_3;
  MG_FA fa_2_55_0(
    .a(pp_2_55_0),
    .b(pp_2_55_1),
    .cin(pp_2_55_2),
    .sum(pp_3_55_0),
    .cout(pp_3_56_0)
  );

  assign pp_3_55_1 = pp_2_55_3;
  assign pp_3_55_2 = pp_2_55_4;
  assign pp_3_56_1 = pp_2_56_0;
  assign pp_3_56_2 = pp_2_56_1;
  assign pp_3_56_3 = pp_2_56_2;
  assign pp_3_56_4 = pp_2_56_3;
  assign pp_3_56_5 = pp_2_56_4;
  MG_FA fa_2_57_0(
    .a(pp_2_57_0),
    .b(pp_2_57_1),
    .cin(pp_2_57_2),
    .sum(pp_3_57_0),
    .cout(pp_3_58_0)
  );

  assign pp_3_57_1 = pp_2_57_3;
  assign pp_3_57_2 = pp_2_57_4;
  MG_FA fa_2_58_0(
    .a(pp_2_58_0),
    .b(pp_2_58_1),
    .cin(pp_2_58_2),
    .sum(pp_3_58_1),
    .cout(pp_3_59_0)
  );

  MG_FA fa_2_59_0(
    .a(pp_2_59_0),
    .b(pp_2_59_1),
    .cin(pp_2_59_2),
    .sum(pp_3_59_1),
    .cout(pp_3_60_0)
  );

  MG_FA fa_2_59_1(
    .a(pp_2_59_3),
    .b(pp_2_59_4),
    .cin(pp_2_59_5),
    .sum(pp_3_59_2),
    .cout(pp_3_60_1)
  );

  assign pp_3_60_2 = pp_2_60_0;
  MG_FA fa_2_61_0(
    .a(pp_2_61_0),
    .b(pp_2_61_1),
    .cin(pp_2_61_2),
    .sum(pp_3_61_0),
    .cout(pp_3_62_0)
  );

  assign pp_3_62_1 = pp_2_62_0;
  assign pp_4_0_0 = pp_3_0_0;
  assign pp_4_1_0 = pp_3_1_0;
  assign pp_4_1_1 = pp_3_1_1;
  assign pp_4_2_0 = pp_3_2_0;
  assign pp_4_2_1 = pp_3_2_1;
  assign pp_4_2_2 = pp_3_2_2;
  MG_FA fa_3_3_0(
    .a(pp_3_3_0),
    .b(pp_3_3_1),
    .cin(pp_3_3_2),
    .sum(pp_4_3_0),
    .cout(pp_4_4_0)
  );

  MG_HA ha_3_4_0(
    .a(pp_3_4_0),
    .b(pp_3_4_1),
    .sum(pp_4_4_1),
    .cout(pp_4_5_0)
  );

  MG_HA ha_3_5_0(
    .a(pp_3_5_0),
    .b(pp_3_5_1),
    .sum(pp_4_5_1),
    .cout(pp_4_6_0)
  );

  MG_FA fa_3_6_0(
    .a(pp_3_6_0),
    .b(pp_3_6_1),
    .cin(pp_3_6_2),
    .sum(pp_4_6_1),
    .cout(pp_4_7_0)
  );

  assign pp_4_6_2 = pp_3_6_3;
  MG_FA fa_3_7_0(
    .a(pp_3_7_0),
    .b(pp_3_7_1),
    .cin(pp_3_7_2),
    .sum(pp_4_7_1),
    .cout(pp_4_8_0)
  );

  assign pp_4_7_2 = pp_3_7_3;
  MG_FA fa_3_8_0(
    .a(pp_3_8_0),
    .b(pp_3_8_1),
    .cin(pp_3_8_2),
    .sum(pp_4_8_1),
    .cout(pp_4_9_0)
  );

  MG_FA fa_3_8_1(
    .a(pp_3_8_3),
    .b(pp_3_8_4),
    .cin(pp_3_8_5),
    .sum(pp_4_8_2),
    .cout(pp_4_9_1)
  );

  MG_FA fa_3_9_0(
    .a(pp_3_9_0),
    .b(pp_3_9_1),
    .cin(pp_3_9_2),
    .sum(pp_4_9_2),
    .cout(pp_4_10_0)
  );

  MG_FA fa_3_10_0(
    .a(pp_3_10_0),
    .b(pp_3_10_1),
    .cin(pp_3_10_2),
    .sum(pp_4_10_1),
    .cout(pp_4_11_0)
  );

  MG_HA ha_3_10_1(
    .a(pp_3_10_3),
    .b(pp_3_10_4),
    .sum(pp_4_10_2),
    .cout(pp_4_11_1)
  );

  MG_FA fa_3_11_0(
    .a(pp_3_11_0),
    .b(pp_3_11_1),
    .cin(pp_3_11_2),
    .sum(pp_4_11_2),
    .cout(pp_4_12_0)
  );

  MG_FA fa_3_11_1(
    .a(pp_3_11_3),
    .b(pp_3_11_4),
    .cin(pp_3_11_5),
    .sum(pp_4_11_3),
    .cout(pp_4_12_1)
  );

  MG_FA fa_3_12_0(
    .a(pp_3_12_0),
    .b(pp_3_12_1),
    .cin(pp_3_12_2),
    .sum(pp_4_12_2),
    .cout(pp_4_13_0)
  );

  MG_FA fa_3_13_0(
    .a(pp_3_13_0),
    .b(pp_3_13_1),
    .cin(pp_3_13_2),
    .sum(pp_4_13_1),
    .cout(pp_4_14_0)
  );

  MG_FA fa_3_14_0(
    .a(pp_3_14_0),
    .b(pp_3_14_1),
    .cin(pp_3_14_2),
    .sum(pp_4_14_1),
    .cout(pp_4_15_0)
  );

  MG_FA fa_3_14_1(
    .a(pp_3_14_3),
    .b(pp_3_14_4),
    .cin(pp_3_14_5),
    .sum(pp_4_14_2),
    .cout(pp_4_15_1)
  );

  MG_FA fa_3_14_2(
    .a(pp_3_14_6),
    .b(pp_3_14_7),
    .cin(pp_3_14_8),
    .sum(pp_4_14_3),
    .cout(pp_4_15_2)
  );

  MG_FA fa_3_15_0(
    .a(pp_3_15_0),
    .b(pp_3_15_1),
    .cin(pp_3_15_2),
    .sum(pp_4_15_3),
    .cout(pp_4_16_0)
  );

  assign pp_4_15_4 = pp_3_15_3;
  assign pp_4_15_5 = pp_3_15_4;
  MG_FA fa_3_16_0(
    .a(pp_3_16_0),
    .b(pp_3_16_1),
    .cin(pp_3_16_2),
    .sum(pp_4_16_1),
    .cout(pp_4_17_0)
  );

  MG_FA fa_3_16_1(
    .a(pp_3_16_3),
    .b(pp_3_16_4),
    .cin(pp_3_16_5),
    .sum(pp_4_16_2),
    .cout(pp_4_17_1)
  );

  MG_FA fa_3_16_2(
    .a(pp_3_16_6),
    .b(pp_3_16_7),
    .cin(pp_3_16_8),
    .sum(pp_4_16_3),
    .cout(pp_4_17_2)
  );

  MG_FA fa_3_17_0(
    .a(pp_3_17_0),
    .b(pp_3_17_1),
    .cin(pp_3_17_2),
    .sum(pp_4_17_3),
    .cout(pp_4_18_0)
  );

  MG_FA fa_3_18_0(
    .a(pp_3_18_0),
    .b(pp_3_18_1),
    .cin(pp_3_18_2),
    .sum(pp_4_18_1),
    .cout(pp_4_19_0)
  );

  MG_FA fa_3_18_1(
    .a(pp_3_18_3),
    .b(pp_3_18_4),
    .cin(pp_3_18_5),
    .sum(pp_4_18_2),
    .cout(pp_4_19_1)
  );

  MG_FA fa_3_18_2(
    .a(pp_3_18_6),
    .b(pp_3_18_7),
    .cin(pp_3_18_8),
    .sum(pp_4_18_3),
    .cout(pp_4_19_2)
  );

  assign pp_4_18_4 = pp_3_18_9;
  assign pp_4_18_5 = pp_3_18_10;
  MG_FA fa_3_19_0(
    .a(pp_3_19_0),
    .b(pp_3_19_1),
    .cin(pp_3_19_2),
    .sum(pp_4_19_3),
    .cout(pp_4_20_0)
  );

  MG_FA fa_3_20_0(
    .a(pp_3_20_0),
    .b(pp_3_20_1),
    .cin(pp_3_20_2),
    .sum(pp_4_20_1),
    .cout(pp_4_21_0)
  );

  MG_FA fa_3_20_1(
    .a(pp_3_20_3),
    .b(pp_3_20_4),
    .cin(pp_3_20_5),
    .sum(pp_4_20_2),
    .cout(pp_4_21_1)
  );

  MG_FA fa_3_21_0(
    .a(pp_3_21_0),
    .b(pp_3_21_1),
    .cin(pp_3_21_2),
    .sum(pp_4_21_2),
    .cout(pp_4_22_0)
  );

  MG_FA fa_3_21_1(
    .a(pp_3_21_3),
    .b(pp_3_21_4),
    .cin(pp_3_21_5),
    .sum(pp_4_21_3),
    .cout(pp_4_22_1)
  );

  MG_FA fa_3_21_2(
    .a(pp_3_21_6),
    .b(pp_3_21_7),
    .cin(pp_3_21_8),
    .sum(pp_4_21_4),
    .cout(pp_4_22_2)
  );

  MG_FA fa_3_22_0(
    .a(pp_3_22_0),
    .b(pp_3_22_1),
    .cin(pp_3_22_2),
    .sum(pp_4_22_3),
    .cout(pp_4_23_0)
  );

  MG_FA fa_3_22_1(
    .a(pp_3_22_3),
    .b(pp_3_22_4),
    .cin(pp_3_22_5),
    .sum(pp_4_22_4),
    .cout(pp_4_23_1)
  );

  MG_FA fa_3_22_2(
    .a(pp_3_22_6),
    .b(pp_3_22_7),
    .cin(pp_3_22_8),
    .sum(pp_4_22_5),
    .cout(pp_4_23_2)
  );

  assign pp_4_22_6 = pp_3_22_9;
  assign pp_4_22_7 = pp_3_22_10;
  MG_FA fa_3_23_0(
    .a(pp_3_23_0),
    .b(pp_3_23_1),
    .cin(pp_3_23_2),
    .sum(pp_4_23_3),
    .cout(pp_4_24_0)
  );

  MG_FA fa_3_23_1(
    .a(pp_3_23_3),
    .b(pp_3_23_4),
    .cin(pp_3_23_5),
    .sum(pp_4_23_4),
    .cout(pp_4_24_1)
  );

  MG_FA fa_3_23_2(
    .a(pp_3_23_6),
    .b(pp_3_23_7),
    .cin(pp_3_23_8),
    .sum(pp_4_23_5),
    .cout(pp_4_24_2)
  );

  MG_FA fa_3_24_0(
    .a(pp_3_24_0),
    .b(pp_3_24_1),
    .cin(pp_3_24_2),
    .sum(pp_4_24_3),
    .cout(pp_4_25_0)
  );

  assign pp_4_24_4 = pp_3_24_3;
  assign pp_4_24_5 = pp_3_24_4;
  MG_FA fa_3_25_0(
    .a(pp_3_25_0),
    .b(pp_3_25_1),
    .cin(pp_3_25_2),
    .sum(pp_4_25_1),
    .cout(pp_4_26_0)
  );

  MG_FA fa_3_25_1(
    .a(pp_3_25_3),
    .b(pp_3_25_4),
    .cin(pp_3_25_5),
    .sum(pp_4_25_2),
    .cout(pp_4_26_1)
  );

  MG_FA fa_3_25_2(
    .a(pp_3_25_6),
    .b(pp_3_25_7),
    .cin(pp_3_25_8),
    .sum(pp_4_25_3),
    .cout(pp_4_26_2)
  );

  MG_FA fa_3_25_3(
    .a(pp_3_25_9),
    .b(pp_3_25_10),
    .cin(pp_3_25_11),
    .sum(pp_4_25_4),
    .cout(pp_4_26_3)
  );

  MG_FA fa_3_25_4(
    .a(pp_3_25_12),
    .b(pp_3_25_13),
    .cin(pp_3_25_14),
    .sum(pp_4_25_5),
    .cout(pp_4_26_4)
  );

  MG_FA fa_3_26_0(
    .a(pp_3_26_0),
    .b(pp_3_26_1),
    .cin(pp_3_26_2),
    .sum(pp_4_26_5),
    .cout(pp_4_27_0)
  );

  MG_FA fa_3_26_1(
    .a(pp_3_26_3),
    .b(pp_3_26_4),
    .cin(pp_3_26_5),
    .sum(pp_4_26_6),
    .cout(pp_4_27_1)
  );

  assign pp_4_26_7 = pp_3_26_6;
  assign pp_4_26_8 = pp_3_26_7;
  MG_FA fa_3_27_0(
    .a(pp_3_27_0),
    .b(pp_3_27_1),
    .cin(pp_3_27_2),
    .sum(pp_4_27_2),
    .cout(pp_4_28_0)
  );

  MG_FA fa_3_27_1(
    .a(pp_3_27_3),
    .b(pp_3_27_4),
    .cin(pp_3_27_5),
    .sum(pp_4_27_3),
    .cout(pp_4_28_1)
  );

  MG_FA fa_3_27_2(
    .a(pp_3_27_6),
    .b(pp_3_27_7),
    .cin(pp_3_27_8),
    .sum(pp_4_27_4),
    .cout(pp_4_28_2)
  );

  MG_FA fa_3_28_0(
    .a(pp_3_28_0),
    .b(pp_3_28_1),
    .cin(pp_3_28_2),
    .sum(pp_4_28_3),
    .cout(pp_4_29_0)
  );

  MG_FA fa_3_28_1(
    .a(pp_3_28_3),
    .b(pp_3_28_4),
    .cin(pp_3_28_5),
    .sum(pp_4_28_4),
    .cout(pp_4_29_1)
  );

  MG_FA fa_3_28_2(
    .a(pp_3_28_6),
    .b(pp_3_28_8),
    .cin(pp_3_28_7),
    .sum(pp_4_28_5),
    .cout(pp_4_29_2)
  );

  MG_FA fa_3_29_0(
    .a(pp_3_29_0),
    .b(pp_3_29_1),
    .cin(pp_3_29_2),
    .sum(pp_4_29_3),
    .cout(pp_4_30_0)
  );

  MG_FA fa_3_29_1(
    .a(pp_3_29_3),
    .b(pp_3_29_4),
    .cin(pp_3_29_5),
    .sum(pp_4_29_4),
    .cout(pp_4_30_1)
  );

  MG_FA fa_3_29_2(
    .a(pp_3_29_6),
    .b(pp_3_29_7),
    .cin(pp_3_29_8),
    .sum(pp_4_29_5),
    .cout(pp_4_30_2)
  );

  MG_FA fa_3_30_0(
    .a(pp_3_30_0),
    .b(pp_3_30_1),
    .cin(pp_3_30_2),
    .sum(pp_4_30_3),
    .cout(pp_4_31_0)
  );

  MG_FA fa_3_30_1(
    .a(pp_3_30_3),
    .b(pp_3_30_4),
    .cin(pp_3_30_5),
    .sum(pp_4_30_4),
    .cout(pp_4_31_1)
  );

  MG_FA fa_3_30_2(
    .a(pp_3_30_6),
    .b(pp_3_30_7),
    .cin(pp_3_30_8),
    .sum(pp_4_30_5),
    .cout(pp_4_31_2)
  );

  MG_FA fa_3_31_0(
    .a(pp_3_31_0),
    .b(pp_3_31_1),
    .cin(pp_3_31_2),
    .sum(pp_4_31_3),
    .cout(pp_4_32_0)
  );

  MG_FA fa_3_31_1(
    .a(pp_3_31_3),
    .b(pp_3_31_4),
    .cin(pp_3_31_5),
    .sum(pp_4_31_4),
    .cout(pp_4_32_1)
  );

  MG_FA fa_3_31_2(
    .a(pp_3_31_6),
    .b(pp_3_31_7),
    .cin(pp_3_31_8),
    .sum(pp_4_31_5),
    .cout(pp_4_32_2)
  );

  MG_FA fa_3_32_0(
    .a(pp_3_32_0),
    .b(pp_3_32_1),
    .cin(pp_3_32_2),
    .sum(pp_4_32_3),
    .cout(pp_4_33_0)
  );

  MG_FA fa_3_32_1(
    .a(pp_3_32_3),
    .b(pp_3_32_4),
    .cin(pp_3_32_5),
    .sum(pp_4_32_4),
    .cout(pp_4_33_1)
  );

  MG_FA fa_3_32_2(
    .a(pp_3_32_6),
    .b(pp_3_32_7),
    .cin(pp_3_32_8),
    .sum(pp_4_32_5),
    .cout(pp_4_33_2)
  );

  assign pp_4_32_6 = pp_3_32_9;
  assign pp_4_32_7 = pp_3_32_10;
  MG_FA fa_3_33_0(
    .a(pp_3_33_0),
    .b(pp_3_33_1),
    .cin(pp_3_33_2),
    .sum(pp_4_33_3),
    .cout(pp_4_34_0)
  );

  MG_FA fa_3_33_1(
    .a(pp_3_33_3),
    .b(pp_3_33_4),
    .cin(pp_3_33_5),
    .sum(pp_4_33_4),
    .cout(pp_4_34_1)
  );

  MG_FA fa_3_33_2(
    .a(pp_3_33_6),
    .b(pp_3_33_7),
    .cin(pp_3_33_8),
    .sum(pp_4_33_5),
    .cout(pp_4_34_2)
  );

  MG_FA fa_3_34_0(
    .a(pp_3_34_0),
    .b(pp_3_34_1),
    .cin(pp_3_34_2),
    .sum(pp_4_34_3),
    .cout(pp_4_35_0)
  );

  MG_FA fa_3_34_1(
    .a(pp_3_34_3),
    .b(pp_3_34_4),
    .cin(pp_3_34_5),
    .sum(pp_4_34_4),
    .cout(pp_4_35_1)
  );

  MG_FA fa_3_34_2(
    .a(pp_3_34_6),
    .b(pp_3_34_7),
    .cin(pp_3_34_8),
    .sum(pp_4_34_5),
    .cout(pp_4_35_2)
  );

  assign pp_4_34_6 = pp_3_34_9;
  MG_FA fa_3_35_0(
    .a(pp_3_35_0),
    .b(pp_3_35_1),
    .cin(pp_3_35_2),
    .sum(pp_4_35_3),
    .cout(pp_4_36_0)
  );

  MG_FA fa_3_35_1(
    .a(pp_3_35_3),
    .b(pp_3_35_4),
    .cin(pp_3_35_5),
    .sum(pp_4_35_4),
    .cout(pp_4_36_1)
  );

  assign pp_4_35_5 = pp_3_35_6;
  assign pp_4_35_6 = pp_3_35_7;
  assign pp_4_35_7 = pp_3_35_8;
  assign pp_4_35_8 = pp_3_35_9;
  MG_FA fa_3_36_0(
    .a(pp_3_36_0),
    .b(pp_3_36_1),
    .cin(pp_3_36_2),
    .sum(pp_4_36_2),
    .cout(pp_4_37_0)
  );

  MG_FA fa_3_36_1(
    .a(pp_3_36_3),
    .b(pp_3_36_4),
    .cin(pp_3_36_5),
    .sum(pp_4_36_3),
    .cout(pp_4_37_1)
  );

  assign pp_4_36_4 = pp_3_36_6;
  assign pp_4_36_5 = pp_3_36_7;
  MG_FA fa_3_37_0(
    .a(pp_3_37_0),
    .b(pp_3_37_1),
    .cin(pp_3_37_2),
    .sum(pp_4_37_2),
    .cout(pp_4_38_0)
  );

  assign pp_4_37_3 = pp_3_37_3;
  assign pp_4_37_4 = pp_3_37_4;
  assign pp_4_37_5 = pp_3_37_5;
  assign pp_4_37_6 = pp_3_37_6;
  assign pp_4_37_7 = pp_3_37_7;
  assign pp_4_37_8 = pp_3_37_8;
  MG_FA fa_3_38_0(
    .a(pp_3_38_0),
    .b(pp_3_38_1),
    .cin(pp_3_38_2),
    .sum(pp_4_38_1),
    .cout(pp_4_39_0)
  );

  MG_FA fa_3_38_1(
    .a(pp_3_38_3),
    .b(pp_3_38_4),
    .cin(pp_3_38_5),
    .sum(pp_4_38_2),
    .cout(pp_4_39_1)
  );

  assign pp_4_38_3 = pp_3_38_6;
  assign pp_4_38_4 = pp_3_38_7;
  assign pp_4_38_5 = pp_3_38_8;
  MG_FA fa_3_39_0(
    .a(pp_3_39_0),
    .b(pp_3_39_1),
    .cin(pp_3_39_2),
    .sum(pp_4_39_2),
    .cout(pp_4_40_0)
  );

  MG_FA fa_3_39_1(
    .a(pp_3_39_3),
    .b(pp_3_39_4),
    .cin(pp_3_39_5),
    .sum(pp_4_39_3),
    .cout(pp_4_40_1)
  );

  MG_FA fa_3_39_2(
    .a(pp_3_39_6),
    .b(pp_3_39_7),
    .cin(pp_3_39_8),
    .sum(pp_4_39_4),
    .cout(pp_4_40_2)
  );

  MG_FA fa_3_40_0(
    .a(pp_3_40_0),
    .b(pp_3_40_1),
    .cin(pp_3_40_2),
    .sum(pp_4_40_3),
    .cout(pp_4_41_0)
  );

  MG_FA fa_3_40_1(
    .a(pp_3_40_3),
    .b(pp_3_40_4),
    .cin(pp_3_40_5),
    .sum(pp_4_40_4),
    .cout(pp_4_41_1)
  );

  assign pp_4_40_5 = pp_3_40_6;
  MG_FA fa_3_41_0(
    .a(pp_3_41_0),
    .b(pp_3_41_1),
    .cin(pp_3_41_2),
    .sum(pp_4_41_2),
    .cout(pp_4_42_0)
  );

  MG_FA fa_3_41_1(
    .a(pp_3_41_3),
    .b(pp_3_41_4),
    .cin(pp_3_41_5),
    .sum(pp_4_41_3),
    .cout(pp_4_42_1)
  );

  MG_FA fa_3_41_2(
    .a(pp_3_41_6),
    .b(pp_3_41_7),
    .cin(pp_3_41_8),
    .sum(pp_4_41_4),
    .cout(pp_4_42_2)
  );

  MG_FA fa_3_41_3(
    .a(pp_3_41_9),
    .b(pp_3_41_10),
    .cin(pp_3_41_11),
    .sum(pp_4_41_5),
    .cout(pp_4_42_3)
  );

  MG_FA fa_3_42_0(
    .a(pp_3_42_0),
    .b(pp_3_42_1),
    .cin(pp_3_42_2),
    .sum(pp_4_42_4),
    .cout(pp_4_43_0)
  );

  assign pp_4_42_5 = pp_3_42_3;
  assign pp_4_42_6 = pp_3_42_4;
  assign pp_4_42_7 = pp_3_42_5;
  MG_FA fa_3_43_0(
    .a(pp_3_43_0),
    .b(pp_3_43_1),
    .cin(pp_3_43_2),
    .sum(pp_4_43_1),
    .cout(pp_4_44_0)
  );

  MG_FA fa_3_43_1(
    .a(pp_3_43_3),
    .b(pp_3_43_4),
    .cin(pp_3_43_5),
    .sum(pp_4_43_2),
    .cout(pp_4_44_1)
  );

  MG_FA fa_3_44_0(
    .a(pp_3_44_0),
    .b(pp_3_44_1),
    .cin(pp_3_44_2),
    .sum(pp_4_44_2),
    .cout(pp_4_45_0)
  );

  MG_FA fa_3_44_1(
    .a(pp_3_44_3),
    .b(pp_3_44_4),
    .cin(pp_3_44_5),
    .sum(pp_4_44_3),
    .cout(pp_4_45_1)
  );

  MG_FA fa_3_44_2(
    .a(pp_3_44_6),
    .b(pp_3_44_7),
    .cin(pp_3_44_8),
    .sum(pp_4_44_4),
    .cout(pp_4_45_2)
  );

  MG_FA fa_3_45_0(
    .a(pp_3_45_0),
    .b(pp_3_45_1),
    .cin(pp_3_45_2),
    .sum(pp_4_45_3),
    .cout(pp_4_46_0)
  );

  MG_FA fa_3_45_1(
    .a(pp_3_45_3),
    .b(pp_3_45_4),
    .cin(pp_3_45_5),
    .sum(pp_4_45_4),
    .cout(pp_4_46_1)
  );

  MG_FA fa_3_45_2(
    .a(pp_3_45_6),
    .b(pp_3_45_7),
    .cin(pp_3_45_8),
    .sum(pp_4_45_5),
    .cout(pp_4_46_2)
  );

  assign pp_4_45_6 = pp_3_45_9;
  MG_FA fa_3_46_0(
    .a(pp_3_46_0),
    .b(pp_3_46_1),
    .cin(pp_3_46_2),
    .sum(pp_4_46_3),
    .cout(pp_4_47_0)
  );

  MG_FA fa_3_46_1(
    .a(pp_3_46_3),
    .b(pp_3_46_4),
    .cin(pp_3_46_5),
    .sum(pp_4_46_4),
    .cout(pp_4_47_1)
  );

  assign pp_4_46_5 = pp_3_46_6;
  assign pp_4_46_6 = pp_3_46_7;
  assign pp_4_46_7 = pp_3_46_8;
  MG_FA fa_3_47_0(
    .a(pp_3_47_0),
    .b(pp_3_47_1),
    .cin(pp_3_47_2),
    .sum(pp_4_47_2),
    .cout(pp_4_48_0)
  );

  MG_FA fa_3_48_0(
    .a(pp_3_48_0),
    .b(pp_3_48_1),
    .cin(pp_3_48_2),
    .sum(pp_4_48_1),
    .cout(pp_4_49_0)
  );

  MG_FA fa_3_48_1(
    .a(pp_3_48_3),
    .b(pp_3_48_4),
    .cin(pp_3_48_5),
    .sum(pp_4_48_2),
    .cout(pp_4_49_1)
  );

  MG_FA fa_3_49_0(
    .a(pp_3_49_0),
    .b(pp_3_49_1),
    .cin(pp_3_49_2),
    .sum(pp_4_49_2),
    .cout(pp_4_50_0)
  );

  MG_FA fa_3_49_1(
    .a(pp_3_49_3),
    .b(pp_3_49_4),
    .cin(pp_3_49_5),
    .sum(pp_4_49_3),
    .cout(pp_4_50_1)
  );

  MG_FA fa_3_50_0(
    .a(pp_3_50_0),
    .b(pp_3_50_1),
    .cin(pp_3_50_2),
    .sum(pp_4_50_2),
    .cout(pp_4_51_0)
  );

  assign pp_4_50_3 = pp_3_50_3;
  assign pp_4_50_4 = pp_3_50_4;
  assign pp_4_50_5 = pp_3_50_5;
  MG_FA fa_3_51_0(
    .a(pp_3_51_0),
    .b(pp_3_51_1),
    .cin(pp_3_51_2),
    .sum(pp_4_51_1),
    .cout(pp_4_52_0)
  );

  MG_FA fa_3_51_1(
    .a(pp_3_51_3),
    .b(pp_3_51_4),
    .cin(pp_3_51_5),
    .sum(pp_4_51_2),
    .cout(pp_4_52_1)
  );

  assign pp_4_52_2 = pp_3_52_0;
  assign pp_4_52_3 = pp_3_52_1;
  assign pp_4_52_4 = pp_3_52_2;
  assign pp_4_52_5 = pp_3_52_3;
  MG_FA fa_3_53_0(
    .a(pp_3_53_0),
    .b(pp_3_53_1),
    .cin(pp_3_53_2),
    .sum(pp_4_53_0),
    .cout(pp_4_54_0)
  );

  MG_FA fa_3_54_0(
    .a(pp_3_54_0),
    .b(pp_3_54_1),
    .cin(pp_3_54_2),
    .sum(pp_4_54_1),
    .cout(pp_4_55_0)
  );

  MG_FA fa_3_54_1(
    .a(pp_3_54_3),
    .b(pp_3_54_4),
    .cin(pp_3_54_5),
    .sum(pp_4_54_2),
    .cout(pp_4_55_1)
  );

  MG_FA fa_3_55_0(
    .a(pp_3_55_0),
    .b(pp_3_55_1),
    .cin(pp_3_55_2),
    .sum(pp_4_55_2),
    .cout(pp_4_56_0)
  );

  MG_FA fa_3_56_0(
    .a(pp_3_56_0),
    .b(pp_3_56_1),
    .cin(pp_3_56_2),
    .sum(pp_4_56_1),
    .cout(pp_4_57_0)
  );

  MG_FA fa_3_56_1(
    .a(pp_3_56_3),
    .b(pp_3_56_4),
    .cin(pp_3_56_5),
    .sum(pp_4_56_2),
    .cout(pp_4_57_1)
  );

  MG_FA fa_3_57_0(
    .a(pp_3_57_0),
    .b(pp_3_57_1),
    .cin(pp_3_57_2),
    .sum(pp_4_57_2),
    .cout(pp_4_58_0)
  );

  assign pp_4_58_1 = pp_3_58_0;
  assign pp_4_58_2 = pp_3_58_1;
  MG_FA fa_3_59_0(
    .a(pp_3_59_0),
    .b(pp_3_59_1),
    .cin(pp_3_59_2),
    .sum(pp_4_59_0),
    .cout(pp_4_60_0)
  );

  MG_FA fa_3_60_0(
    .a(pp_3_60_0),
    .b(pp_3_60_1),
    .cin(pp_3_60_2),
    .sum(pp_4_60_1),
    .cout(pp_4_61_0)
  );

  assign pp_4_61_1 = pp_3_61_0;
  assign pp_4_62_0 = pp_3_62_0;
  assign pp_4_62_1 = pp_3_62_1;
  assign pp_5_0_0 = pp_4_0_0;
  assign pp_5_1_0 = pp_4_1_0;
  assign pp_5_1_1 = pp_4_1_1;
  MG_HA ha_4_2_0(
    .a(pp_4_2_0),
    .b(pp_4_2_1),
    .sum(pp_5_2_0),
    .cout(pp_5_3_0)
  );

  assign pp_5_2_1 = pp_4_2_2;
  assign pp_5_3_1 = pp_4_3_0;
  assign pp_5_4_0 = pp_4_4_0;
  assign pp_5_4_1 = pp_4_4_1;
  assign pp_5_5_0 = pp_4_5_0;
  assign pp_5_5_1 = pp_4_5_1;
  assign pp_5_6_0 = pp_4_6_0;
  assign pp_5_6_1 = pp_4_6_1;
  assign pp_5_6_2 = pp_4_6_2;
  MG_FA fa_4_7_0(
    .a(pp_4_7_0),
    .b(pp_4_7_1),
    .cin(pp_4_7_2),
    .sum(pp_5_7_0),
    .cout(pp_5_8_0)
  );

  MG_FA fa_4_8_0(
    .a(pp_4_8_0),
    .b(pp_4_8_1),
    .cin(pp_4_8_2),
    .sum(pp_5_8_1),
    .cout(pp_5_9_0)
  );

  MG_FA fa_4_9_0(
    .a(pp_4_9_0),
    .b(pp_4_9_1),
    .cin(pp_4_9_2),
    .sum(pp_5_9_1),
    .cout(pp_5_10_0)
  );

  MG_FA fa_4_10_0(
    .a(pp_4_10_0),
    .b(pp_4_10_1),
    .cin(pp_4_10_2),
    .sum(pp_5_10_1),
    .cout(pp_5_11_0)
  );

  MG_HA ha_4_11_0(
    .a(pp_4_11_0),
    .b(pp_4_11_1),
    .sum(pp_5_11_1),
    .cout(pp_5_12_0)
  );

  assign pp_5_11_2 = pp_4_11_2;
  assign pp_5_11_3 = pp_4_11_3;
  MG_FA fa_4_12_0(
    .a(pp_4_12_0),
    .b(pp_4_12_1),
    .cin(pp_4_12_2),
    .sum(pp_5_12_1),
    .cout(pp_5_13_0)
  );

  assign pp_5_13_1 = pp_4_13_0;
  assign pp_5_13_2 = pp_4_13_1;
  MG_FA fa_4_14_0(
    .a(pp_4_14_0),
    .b(pp_4_14_1),
    .cin(pp_4_14_2),
    .sum(pp_5_14_0),
    .cout(pp_5_15_0)
  );

  assign pp_5_14_1 = pp_4_14_3;
  MG_FA fa_4_15_0(
    .a(pp_4_15_0),
    .b(pp_4_15_1),
    .cin(pp_4_15_2),
    .sum(pp_5_15_1),
    .cout(pp_5_16_0)
  );

  MG_FA fa_4_15_1(
    .a(pp_4_15_3),
    .b(pp_4_15_4),
    .cin(pp_4_15_5),
    .sum(pp_5_15_2),
    .cout(pp_5_16_1)
  );

  assign pp_5_16_2 = pp_4_16_0;
  assign pp_5_16_3 = pp_4_16_1;
  assign pp_5_16_4 = pp_4_16_2;
  assign pp_5_16_5 = pp_4_16_3;
  MG_FA fa_4_17_0(
    .a(pp_4_17_0),
    .b(pp_4_17_1),
    .cin(pp_4_17_2),
    .sum(pp_5_17_0),
    .cout(pp_5_18_0)
  );

  assign pp_5_17_1 = pp_4_17_3;
  MG_FA fa_4_18_0(
    .a(pp_4_18_0),
    .b(pp_4_18_1),
    .cin(pp_4_18_2),
    .sum(pp_5_18_1),
    .cout(pp_5_19_0)
  );

  MG_FA fa_4_18_1(
    .a(pp_4_18_3),
    .b(pp_4_18_4),
    .cin(pp_4_18_5),
    .sum(pp_5_18_2),
    .cout(pp_5_19_1)
  );

  assign pp_5_19_2 = pp_4_19_0;
  assign pp_5_19_3 = pp_4_19_1;
  assign pp_5_19_4 = pp_4_19_2;
  assign pp_5_19_5 = pp_4_19_3;
  MG_FA fa_4_20_0(
    .a(pp_4_20_0),
    .b(pp_4_20_1),
    .cin(pp_4_20_2),
    .sum(pp_5_20_0),
    .cout(pp_5_21_0)
  );

  MG_FA fa_4_21_0(
    .a(pp_4_21_0),
    .b(pp_4_21_1),
    .cin(pp_4_21_2),
    .sum(pp_5_21_1),
    .cout(pp_5_22_0)
  );

  MG_HA ha_4_21_1(
    .a(pp_4_21_3),
    .b(pp_4_21_4),
    .sum(pp_5_21_2),
    .cout(pp_5_22_1)
  );

  MG_FA fa_4_22_0(
    .a(pp_4_22_0),
    .b(pp_4_22_1),
    .cin(pp_4_22_2),
    .sum(pp_5_22_2),
    .cout(pp_5_23_0)
  );

  MG_FA fa_4_22_1(
    .a(pp_4_22_3),
    .b(pp_4_22_4),
    .cin(pp_4_22_5),
    .sum(pp_5_22_3),
    .cout(pp_5_23_1)
  );

  assign pp_5_22_4 = pp_4_22_6;
  assign pp_5_22_5 = pp_4_22_7;
  MG_FA fa_4_23_0(
    .a(pp_4_23_0),
    .b(pp_4_23_1),
    .cin(pp_4_23_2),
    .sum(pp_5_23_2),
    .cout(pp_5_24_0)
  );

  MG_FA fa_4_23_1(
    .a(pp_4_23_3),
    .b(pp_4_23_4),
    .cin(pp_4_23_5),
    .sum(pp_5_23_3),
    .cout(pp_5_24_1)
  );

  MG_FA fa_4_24_0(
    .a(pp_4_24_0),
    .b(pp_4_24_1),
    .cin(pp_4_24_2),
    .sum(pp_5_24_2),
    .cout(pp_5_25_0)
  );

  MG_FA fa_4_24_1(
    .a(pp_4_24_3),
    .b(pp_4_24_4),
    .cin(pp_4_24_5),
    .sum(pp_5_24_3),
    .cout(pp_5_25_1)
  );

  MG_FA fa_4_25_0(
    .a(pp_4_25_0),
    .b(pp_4_25_1),
    .cin(pp_4_25_2),
    .sum(pp_5_25_2),
    .cout(pp_5_26_0)
  );

  MG_FA fa_4_25_1(
    .a(pp_4_25_3),
    .b(pp_4_25_4),
    .cin(pp_4_25_5),
    .sum(pp_5_25_3),
    .cout(pp_5_26_1)
  );

  MG_FA fa_4_26_0(
    .a(pp_4_26_0),
    .b(pp_4_26_1),
    .cin(pp_4_26_2),
    .sum(pp_5_26_2),
    .cout(pp_5_27_0)
  );

  assign pp_5_26_3 = pp_4_26_3;
  assign pp_5_26_4 = pp_4_26_4;
  assign pp_5_26_5 = pp_4_26_5;
  assign pp_5_26_6 = pp_4_26_6;
  assign pp_5_26_7 = pp_4_26_7;
  assign pp_5_26_8 = pp_4_26_8;
  MG_FA fa_4_27_0(
    .a(pp_4_27_0),
    .b(pp_4_27_1),
    .cin(pp_4_27_2),
    .sum(pp_5_27_1),
    .cout(pp_5_28_0)
  );

  assign pp_5_27_2 = pp_4_27_3;
  assign pp_5_27_3 = pp_4_27_4;
  MG_FA fa_4_28_0(
    .a(pp_4_28_0),
    .b(pp_4_28_1),
    .cin(pp_4_28_2),
    .sum(pp_5_28_1),
    .cout(pp_5_29_0)
  );

  MG_FA fa_4_28_1(
    .a(pp_4_28_3),
    .b(pp_4_28_4),
    .cin(pp_4_28_5),
    .sum(pp_5_28_2),
    .cout(pp_5_29_1)
  );

  MG_FA fa_4_29_0(
    .a(pp_4_29_0),
    .b(pp_4_29_1),
    .cin(pp_4_29_2),
    .sum(pp_5_29_2),
    .cout(pp_5_30_0)
  );

  MG_HA ha_4_29_1(
    .a(pp_4_29_3),
    .b(pp_4_29_4),
    .sum(pp_5_29_3),
    .cout(pp_5_30_1)
  );

  assign pp_5_29_4 = pp_4_29_5;
  MG_FA fa_4_30_0(
    .a(pp_4_30_0),
    .b(pp_4_30_1),
    .cin(pp_4_30_2),
    .sum(pp_5_30_2),
    .cout(pp_5_31_0)
  );

  MG_FA fa_4_30_1(
    .a(pp_4_30_3),
    .b(pp_4_30_4),
    .cin(pp_4_30_5),
    .sum(pp_5_30_3),
    .cout(pp_5_31_1)
  );

  MG_FA fa_4_31_0(
    .a(pp_4_31_0),
    .b(pp_4_31_1),
    .cin(pp_4_31_2),
    .sum(pp_5_31_2),
    .cout(pp_5_32_0)
  );

  assign pp_5_31_3 = pp_4_31_3;
  assign pp_5_31_4 = pp_4_31_4;
  assign pp_5_31_5 = pp_4_31_5;
  MG_FA fa_4_32_0(
    .a(pp_4_32_0),
    .b(pp_4_32_1),
    .cin(pp_4_32_2),
    .sum(pp_5_32_1),
    .cout(pp_5_33_0)
  );

  MG_FA fa_4_32_1(
    .a(pp_4_32_3),
    .b(pp_4_32_4),
    .cin(pp_4_32_5),
    .sum(pp_5_32_2),
    .cout(pp_5_33_1)
  );

  assign pp_5_32_3 = pp_4_32_6;
  assign pp_5_32_4 = pp_4_32_7;
  MG_FA fa_4_33_0(
    .a(pp_4_33_0),
    .b(pp_4_33_1),
    .cin(pp_4_33_2),
    .sum(pp_5_33_2),
    .cout(pp_5_34_0)
  );

  MG_FA fa_4_33_1(
    .a(pp_4_33_3),
    .b(pp_4_33_4),
    .cin(pp_4_33_5),
    .sum(pp_5_33_3),
    .cout(pp_5_34_1)
  );

  assign pp_5_34_2 = pp_4_34_0;
  assign pp_5_34_3 = pp_4_34_1;
  assign pp_5_34_4 = pp_4_34_2;
  assign pp_5_34_5 = pp_4_34_3;
  assign pp_5_34_6 = pp_4_34_4;
  assign pp_5_34_7 = pp_4_34_5;
  assign pp_5_34_8 = pp_4_34_6;
  MG_FA fa_4_35_0(
    .a(pp_4_35_0),
    .b(pp_4_35_1),
    .cin(pp_4_35_2),
    .sum(pp_5_35_0),
    .cout(pp_5_36_0)
  );

  MG_FA fa_4_35_1(
    .a(pp_4_35_3),
    .b(pp_4_35_4),
    .cin(pp_4_35_5),
    .sum(pp_5_35_1),
    .cout(pp_5_36_1)
  );

  MG_FA fa_4_35_2(
    .a(pp_4_35_6),
    .b(pp_4_35_7),
    .cin(pp_4_35_8),
    .sum(pp_5_35_2),
    .cout(pp_5_36_2)
  );

  assign pp_5_36_3 = pp_4_36_0;
  assign pp_5_36_4 = pp_4_36_1;
  assign pp_5_36_5 = pp_4_36_2;
  assign pp_5_36_6 = pp_4_36_3;
  assign pp_5_36_7 = pp_4_36_4;
  assign pp_5_36_8 = pp_4_36_5;
  MG_FA fa_4_37_0(
    .a(pp_4_37_0),
    .b(pp_4_37_1),
    .cin(pp_4_37_2),
    .sum(pp_5_37_0),
    .cout(pp_5_38_0)
  );

  MG_FA fa_4_37_1(
    .a(pp_4_37_3),
    .b(pp_4_37_4),
    .cin(pp_4_37_5),
    .sum(pp_5_37_1),
    .cout(pp_5_38_1)
  );

  MG_FA fa_4_37_2(
    .a(pp_4_37_6),
    .b(pp_4_37_7),
    .cin(pp_4_37_8),
    .sum(pp_5_37_2),
    .cout(pp_5_38_2)
  );

  assign pp_5_38_3 = pp_4_38_0;
  assign pp_5_38_4 = pp_4_38_1;
  assign pp_5_38_5 = pp_4_38_2;
  assign pp_5_38_6 = pp_4_38_3;
  assign pp_5_38_7 = pp_4_38_4;
  assign pp_5_38_8 = pp_4_38_5;
  MG_FA fa_4_39_0(
    .a(pp_4_39_0),
    .b(pp_4_39_1),
    .cin(pp_4_39_2),
    .sum(pp_5_39_0),
    .cout(pp_5_40_0)
  );

  assign pp_5_39_1 = pp_4_39_3;
  assign pp_5_39_2 = pp_4_39_4;
  MG_FA fa_4_40_0(
    .a(pp_4_40_0),
    .b(pp_4_40_1),
    .cin(pp_4_40_2),
    .sum(pp_5_40_1),
    .cout(pp_5_41_0)
  );

  MG_FA fa_4_40_1(
    .a(pp_4_40_3),
    .b(pp_4_40_4),
    .cin(pp_4_40_5),
    .sum(pp_5_40_2),
    .cout(pp_5_41_1)
  );

  assign pp_5_41_2 = pp_4_41_0;
  assign pp_5_41_3 = pp_4_41_1;
  assign pp_5_41_4 = pp_4_41_2;
  assign pp_5_41_5 = pp_4_41_3;
  assign pp_5_41_6 = pp_4_41_4;
  assign pp_5_41_7 = pp_4_41_5;
  MG_FA fa_4_42_0(
    .a(pp_4_42_0),
    .b(pp_4_42_1),
    .cin(pp_4_42_2),
    .sum(pp_5_42_0),
    .cout(pp_5_43_0)
  );

  MG_FA fa_4_42_1(
    .a(pp_4_42_3),
    .b(pp_4_42_4),
    .cin(pp_4_42_5),
    .sum(pp_5_42_1),
    .cout(pp_5_43_1)
  );

  assign pp_5_42_2 = pp_4_42_6;
  assign pp_5_42_3 = pp_4_42_7;
  MG_FA fa_4_43_0(
    .a(pp_4_43_0),
    .b(pp_4_43_1),
    .cin(pp_4_43_2),
    .sum(pp_5_43_2),
    .cout(pp_5_44_0)
  );

  assign pp_5_44_1 = pp_4_44_0;
  assign pp_5_44_2 = pp_4_44_1;
  assign pp_5_44_3 = pp_4_44_2;
  assign pp_5_44_4 = pp_4_44_3;
  assign pp_5_44_5 = pp_4_44_4;
  MG_FA fa_4_45_0(
    .a(pp_4_45_0),
    .b(pp_4_45_1),
    .cin(pp_4_45_2),
    .sum(pp_5_45_0),
    .cout(pp_5_46_0)
  );

  MG_FA fa_4_45_1(
    .a(pp_4_45_3),
    .b(pp_4_45_4),
    .cin(pp_4_45_5),
    .sum(pp_5_45_1),
    .cout(pp_5_46_1)
  );

  assign pp_5_45_2 = pp_4_45_6;
  MG_FA fa_4_46_0(
    .a(pp_4_46_0),
    .b(pp_4_46_1),
    .cin(pp_4_46_2),
    .sum(pp_5_46_2),
    .cout(pp_5_47_0)
  );

  MG_FA fa_4_46_1(
    .a(pp_4_46_3),
    .b(pp_4_46_4),
    .cin(pp_4_46_5),
    .sum(pp_5_46_3),
    .cout(pp_5_47_1)
  );

  assign pp_5_46_4 = pp_4_46_6;
  assign pp_5_46_5 = pp_4_46_7;
  MG_FA fa_4_47_0(
    .a(pp_4_47_0),
    .b(pp_4_47_1),
    .cin(pp_4_47_2),
    .sum(pp_5_47_2),
    .cout(pp_5_48_0)
  );

  assign pp_5_48_1 = pp_4_48_0;
  assign pp_5_48_2 = pp_4_48_1;
  assign pp_5_48_3 = pp_4_48_2;
  MG_FA fa_4_49_0(
    .a(pp_4_49_0),
    .b(pp_4_49_1),
    .cin(pp_4_49_2),
    .sum(pp_5_49_0),
    .cout(pp_5_50_0)
  );

  assign pp_5_49_1 = pp_4_49_3;
  assign pp_5_50_1 = pp_4_50_0;
  assign pp_5_50_2 = pp_4_50_1;
  assign pp_5_50_3 = pp_4_50_2;
  assign pp_5_50_4 = pp_4_50_3;
  assign pp_5_50_5 = pp_4_50_4;
  assign pp_5_50_6 = pp_4_50_5;
  MG_FA fa_4_51_0(
    .a(pp_4_51_0),
    .b(pp_4_51_1),
    .cin(pp_4_51_2),
    .sum(pp_5_51_0),
    .cout(pp_5_52_0)
  );

  assign pp_5_52_1 = pp_4_52_0;
  assign pp_5_52_2 = pp_4_52_1;
  assign pp_5_52_3 = pp_4_52_2;
  assign pp_5_52_4 = pp_4_52_3;
  assign pp_5_52_5 = pp_4_52_4;
  assign pp_5_52_6 = pp_4_52_5;
  assign pp_5_53_0 = pp_4_53_0;
  assign pp_5_54_0 = pp_4_54_0;
  assign pp_5_54_1 = pp_4_54_1;
  assign pp_5_54_2 = pp_4_54_2;
  assign pp_5_55_0 = pp_4_55_0;
  assign pp_5_55_1 = pp_4_55_1;
  assign pp_5_55_2 = pp_4_55_2;
  assign pp_5_56_0 = pp_4_56_0;
  assign pp_5_56_1 = pp_4_56_1;
  assign pp_5_56_2 = pp_4_56_2;
  MG_FA fa_4_57_0(
    .a(pp_4_57_0),
    .b(pp_4_57_1),
    .cin(pp_4_57_2),
    .sum(pp_5_57_0),
    .cout(pp_5_58_0)
  );

  MG_FA fa_4_58_0(
    .a(pp_4_58_0),
    .b(pp_4_58_1),
    .cin(pp_4_58_2),
    .sum(pp_5_58_1),
    .cout(pp_5_59_0)
  );

  assign pp_5_59_1 = pp_4_59_0;
  assign pp_5_60_0 = pp_4_60_0;
  assign pp_5_60_1 = pp_4_60_1;
  assign pp_5_61_0 = pp_4_61_0;
  assign pp_5_61_1 = pp_4_61_1;
  assign pp_5_62_0 = pp_4_62_0;
  assign pp_5_62_1 = pp_4_62_1;
  assign pp_6_0_0 = pp_5_0_0;
  assign pp_6_1_0 = pp_5_1_0;
  assign pp_6_1_1 = pp_5_1_1;
  assign pp_6_2_0 = pp_5_2_0;
  assign pp_6_2_1 = pp_5_2_1;
  assign pp_6_3_0 = pp_5_3_0;
  assign pp_6_3_1 = pp_5_3_1;
  assign pp_6_4_0 = pp_5_4_0;
  assign pp_6_4_1 = pp_5_4_1;
  assign pp_6_5_0 = pp_5_5_0;
  assign pp_6_5_1 = pp_5_5_1;
  assign pp_6_6_0 = pp_5_6_0;
  assign pp_6_6_1 = pp_5_6_1;
  assign pp_6_6_2 = pp_5_6_2;
  assign pp_6_7_0 = pp_5_7_0;
  assign pp_6_8_0 = pp_5_8_0;
  assign pp_6_8_1 = pp_5_8_1;
  assign pp_6_9_0 = pp_5_9_0;
  assign pp_6_9_1 = pp_5_9_1;
  assign pp_6_10_0 = pp_5_10_0;
  assign pp_6_10_1 = pp_5_10_1;
  assign pp_6_11_0 = pp_5_11_0;
  assign pp_6_11_1 = pp_5_11_1;
  assign pp_6_11_2 = pp_5_11_2;
  assign pp_6_11_3 = pp_5_11_3;
  MG_HA ha_5_12_0(
    .a(pp_5_12_0),
    .b(pp_5_12_1),
    .sum(pp_6_12_0),
    .cout(pp_6_13_0)
  );

  MG_FA fa_5_13_0(
    .a(pp_5_13_0),
    .b(pp_5_13_1),
    .cin(pp_5_13_2),
    .sum(pp_6_13_1),
    .cout(pp_6_14_0)
  );

  assign pp_6_14_1 = pp_5_14_0;
  assign pp_6_14_2 = pp_5_14_1;
  MG_FA fa_5_15_0(
    .a(pp_5_15_0),
    .b(pp_5_15_1),
    .cin(pp_5_15_2),
    .sum(pp_6_15_0),
    .cout(pp_6_16_0)
  );

  MG_FA fa_5_16_0(
    .a(pp_5_16_0),
    .b(pp_5_16_1),
    .cin(pp_5_16_2),
    .sum(pp_6_16_1),
    .cout(pp_6_17_0)
  );

  MG_FA fa_5_16_1(
    .a(pp_5_16_3),
    .b(pp_5_16_4),
    .cin(pp_5_16_5),
    .sum(pp_6_16_2),
    .cout(pp_6_17_1)
  );

  MG_HA ha_5_17_0(
    .a(pp_5_17_0),
    .b(pp_5_17_1),
    .sum(pp_6_17_2),
    .cout(pp_6_18_0)
  );

  MG_FA fa_5_18_0(
    .a(pp_5_18_0),
    .b(pp_5_18_1),
    .cin(pp_5_18_2),
    .sum(pp_6_18_1),
    .cout(pp_6_19_0)
  );

  MG_FA fa_5_19_0(
    .a(pp_5_19_0),
    .b(pp_5_19_1),
    .cin(pp_5_19_2),
    .sum(pp_6_19_1),
    .cout(pp_6_20_0)
  );

  MG_FA fa_5_19_1(
    .a(pp_5_19_3),
    .b(pp_5_19_4),
    .cin(pp_5_19_5),
    .sum(pp_6_19_2),
    .cout(pp_6_20_1)
  );

  assign pp_6_20_2 = pp_5_20_0;
  assign pp_6_21_0 = pp_5_21_0;
  assign pp_6_21_1 = pp_5_21_1;
  assign pp_6_21_2 = pp_5_21_2;
  MG_FA fa_5_22_0(
    .a(pp_5_22_0),
    .b(pp_5_22_1),
    .cin(pp_5_22_2),
    .sum(pp_6_22_0),
    .cout(pp_6_23_0)
  );

  MG_FA fa_5_22_1(
    .a(pp_5_22_3),
    .b(pp_5_22_4),
    .cin(pp_5_22_5),
    .sum(pp_6_22_1),
    .cout(pp_6_23_1)
  );

  MG_FA fa_5_23_0(
    .a(pp_5_23_0),
    .b(pp_5_23_1),
    .cin(pp_5_23_2),
    .sum(pp_6_23_2),
    .cout(pp_6_24_0)
  );

  assign pp_6_23_3 = pp_5_23_3;
  MG_FA fa_5_24_0(
    .a(pp_5_24_0),
    .b(pp_5_24_1),
    .cin(pp_5_24_2),
    .sum(pp_6_24_1),
    .cout(pp_6_25_0)
  );

  assign pp_6_24_2 = pp_5_24_3;
  MG_HA ha_5_25_0(
    .a(pp_5_25_0),
    .b(pp_5_25_1),
    .sum(pp_6_25_1),
    .cout(pp_6_26_0)
  );

  assign pp_6_25_2 = pp_5_25_2;
  assign pp_6_25_3 = pp_5_25_3;
  MG_FA fa_5_26_0(
    .a(pp_5_26_0),
    .b(pp_5_26_1),
    .cin(pp_5_26_2),
    .sum(pp_6_26_1),
    .cout(pp_6_27_0)
  );

  MG_FA fa_5_26_1(
    .a(pp_5_26_3),
    .b(pp_5_26_4),
    .cin(pp_5_26_5),
    .sum(pp_6_26_2),
    .cout(pp_6_27_1)
  );

  MG_FA fa_5_26_2(
    .a(pp_5_26_6),
    .b(pp_5_26_7),
    .cin(pp_5_26_8),
    .sum(pp_6_26_3),
    .cout(pp_6_27_2)
  );

  MG_FA fa_5_27_0(
    .a(pp_5_27_0),
    .b(pp_5_27_1),
    .cin(pp_5_27_2),
    .sum(pp_6_27_3),
    .cout(pp_6_28_0)
  );

  assign pp_6_27_4 = pp_5_27_3;
  MG_FA fa_5_28_0(
    .a(pp_5_28_0),
    .b(pp_5_28_1),
    .cin(pp_5_28_2),
    .sum(pp_6_28_1),
    .cout(pp_6_29_0)
  );

  MG_FA fa_5_29_0(
    .a(pp_5_29_0),
    .b(pp_5_29_1),
    .cin(pp_5_29_2),
    .sum(pp_6_29_1),
    .cout(pp_6_30_0)
  );

  assign pp_6_29_2 = pp_5_29_3;
  assign pp_6_29_3 = pp_5_29_4;
  MG_FA fa_5_30_0(
    .a(pp_5_30_0),
    .b(pp_5_30_1),
    .cin(pp_5_30_2),
    .sum(pp_6_30_1),
    .cout(pp_6_31_0)
  );

  assign pp_6_30_2 = pp_5_30_3;
  MG_FA fa_5_31_0(
    .a(pp_5_31_0),
    .b(pp_5_31_1),
    .cin(pp_5_31_2),
    .sum(pp_6_31_1),
    .cout(pp_6_32_0)
  );

  MG_FA fa_5_31_1(
    .a(pp_5_31_3),
    .b(pp_5_31_4),
    .cin(pp_5_31_5),
    .sum(pp_6_31_2),
    .cout(pp_6_32_1)
  );

  MG_FA fa_5_32_0(
    .a(pp_5_32_0),
    .b(pp_5_32_1),
    .cin(pp_5_32_2),
    .sum(pp_6_32_2),
    .cout(pp_6_33_0)
  );

  assign pp_6_32_3 = pp_5_32_3;
  assign pp_6_32_4 = pp_5_32_4;
  MG_FA fa_5_33_0(
    .a(pp_5_33_0),
    .b(pp_5_33_1),
    .cin(pp_5_33_2),
    .sum(pp_6_33_1),
    .cout(pp_6_34_0)
  );

  assign pp_6_33_2 = pp_5_33_3;
  MG_FA fa_5_34_0(
    .a(pp_5_34_0),
    .b(pp_5_34_2),
    .cin(pp_5_34_1),
    .sum(pp_6_34_1),
    .cout(pp_6_35_0)
  );

  MG_FA fa_5_34_1(
    .a(pp_5_34_3),
    .b(pp_5_34_4),
    .cin(pp_5_34_5),
    .sum(pp_6_34_2),
    .cout(pp_6_35_1)
  );

  MG_FA fa_5_34_2(
    .a(pp_5_34_6),
    .b(pp_5_34_7),
    .cin(pp_5_34_8),
    .sum(pp_6_34_3),
    .cout(pp_6_35_2)
  );

  MG_FA fa_5_35_0(
    .a(pp_5_35_0),
    .b(pp_5_35_1),
    .cin(pp_5_35_2),
    .sum(pp_6_35_3),
    .cout(pp_6_36_0)
  );

  MG_FA fa_5_36_0(
    .a(pp_5_36_0),
    .b(pp_5_36_1),
    .cin(pp_5_36_2),
    .sum(pp_6_36_1),
    .cout(pp_6_37_0)
  );

  MG_FA fa_5_36_1(
    .a(pp_5_36_3),
    .b(pp_5_36_4),
    .cin(pp_5_36_5),
    .sum(pp_6_36_2),
    .cout(pp_6_37_1)
  );

  MG_FA fa_5_36_2(
    .a(pp_5_36_6),
    .b(pp_5_36_7),
    .cin(pp_5_36_8),
    .sum(pp_6_36_3),
    .cout(pp_6_37_2)
  );

  MG_FA fa_5_37_0(
    .a(pp_5_37_0),
    .b(pp_5_37_1),
    .cin(pp_5_37_2),
    .sum(pp_6_37_3),
    .cout(pp_6_38_0)
  );

  MG_FA fa_5_38_0(
    .a(pp_5_38_0),
    .b(pp_5_38_1),
    .cin(pp_5_38_2),
    .sum(pp_6_38_1),
    .cout(pp_6_39_0)
  );

  MG_FA fa_5_38_1(
    .a(pp_5_38_3),
    .b(pp_5_38_4),
    .cin(pp_5_38_5),
    .sum(pp_6_38_2),
    .cout(pp_6_39_1)
  );

  MG_FA fa_5_38_2(
    .a(pp_5_38_6),
    .b(pp_5_38_7),
    .cin(pp_5_38_8),
    .sum(pp_6_38_3),
    .cout(pp_6_39_2)
  );

  MG_FA fa_5_39_0(
    .a(pp_5_39_0),
    .b(pp_5_39_1),
    .cin(pp_5_39_2),
    .sum(pp_6_39_3),
    .cout(pp_6_40_0)
  );

  MG_FA fa_5_40_0(
    .a(pp_5_40_0),
    .b(pp_5_40_1),
    .cin(pp_5_40_2),
    .sum(pp_6_40_1),
    .cout(pp_6_41_0)
  );

  MG_FA fa_5_41_0(
    .a(pp_5_41_0),
    .b(pp_5_41_1),
    .cin(pp_5_41_2),
    .sum(pp_6_41_1),
    .cout(pp_6_42_0)
  );

  assign pp_6_41_2 = pp_5_41_3;
  assign pp_6_41_3 = pp_5_41_4;
  assign pp_6_41_4 = pp_5_41_5;
  assign pp_6_41_5 = pp_5_41_6;
  assign pp_6_41_6 = pp_5_41_7;
  MG_FA fa_5_42_0(
    .a(pp_5_42_0),
    .b(pp_5_42_1),
    .cin(pp_5_42_2),
    .sum(pp_6_42_1),
    .cout(pp_6_43_0)
  );

  assign pp_6_42_2 = pp_5_42_3;
  MG_FA fa_5_43_0(
    .a(pp_5_43_0),
    .b(pp_5_43_1),
    .cin(pp_5_43_2),
    .sum(pp_6_43_1),
    .cout(pp_6_44_0)
  );

  MG_FA fa_5_44_0(
    .a(pp_5_44_0),
    .b(pp_5_44_1),
    .cin(pp_5_44_2),
    .sum(pp_6_44_1),
    .cout(pp_6_45_0)
  );

  MG_FA fa_5_44_1(
    .a(pp_5_44_3),
    .b(pp_5_44_4),
    .cin(pp_5_44_5),
    .sum(pp_6_44_2),
    .cout(pp_6_45_1)
  );

  assign pp_6_45_2 = pp_5_45_0;
  assign pp_6_45_3 = pp_5_45_1;
  assign pp_6_45_4 = pp_5_45_2;
  MG_FA fa_5_46_0(
    .a(pp_5_46_0),
    .b(pp_5_46_1),
    .cin(pp_5_46_2),
    .sum(pp_6_46_0),
    .cout(pp_6_47_0)
  );

  MG_FA fa_5_46_1(
    .a(pp_5_46_3),
    .b(pp_5_46_4),
    .cin(pp_5_46_5),
    .sum(pp_6_46_1),
    .cout(pp_6_47_1)
  );

  MG_FA fa_5_47_0(
    .a(pp_5_47_0),
    .b(pp_5_47_1),
    .cin(pp_5_47_2),
    .sum(pp_6_47_2),
    .cout(pp_6_48_0)
  );

  MG_FA fa_5_48_0(
    .a(pp_5_48_0),
    .b(pp_5_48_1),
    .cin(pp_5_48_2),
    .sum(pp_6_48_1),
    .cout(pp_6_49_0)
  );

  assign pp_6_48_2 = pp_5_48_3;
  assign pp_6_49_1 = pp_5_49_0;
  assign pp_6_49_2 = pp_5_49_1;
  MG_FA fa_5_50_0(
    .a(pp_5_50_0),
    .b(pp_5_50_1),
    .cin(pp_5_50_2),
    .sum(pp_6_50_0),
    .cout(pp_6_51_0)
  );

  MG_FA fa_5_50_1(
    .a(pp_5_50_3),
    .b(pp_5_50_4),
    .cin(pp_5_50_5),
    .sum(pp_6_50_1),
    .cout(pp_6_51_1)
  );

  assign pp_6_50_2 = pp_5_50_6;
  assign pp_6_51_2 = pp_5_51_0;
  MG_FA fa_5_52_0(
    .a(pp_5_52_0),
    .b(pp_5_52_1),
    .cin(pp_5_52_2),
    .sum(pp_6_52_0),
    .cout(pp_6_53_0)
  );

  MG_FA fa_5_52_1(
    .a(pp_5_52_3),
    .b(pp_5_52_4),
    .cin(pp_5_52_5),
    .sum(pp_6_52_1),
    .cout(pp_6_53_1)
  );

  assign pp_6_52_2 = pp_5_52_6;
  assign pp_6_53_2 = pp_5_53_0;
  MG_FA fa_5_54_0(
    .a(pp_5_54_0),
    .b(pp_5_54_1),
    .cin(pp_5_54_2),
    .sum(pp_6_54_0),
    .cout(pp_6_55_0)
  );

  MG_FA fa_5_55_0(
    .a(pp_5_55_0),
    .b(pp_5_55_1),
    .cin(pp_5_55_2),
    .sum(pp_6_55_1),
    .cout(pp_6_56_0)
  );

  MG_FA fa_5_56_0(
    .a(pp_5_56_0),
    .b(pp_5_56_1),
    .cin(pp_5_56_2),
    .sum(pp_6_56_1),
    .cout(pp_6_57_0)
  );

  assign pp_6_57_1 = pp_5_57_0;
  assign pp_6_58_0 = pp_5_58_0;
  assign pp_6_58_1 = pp_5_58_1;
  assign pp_6_59_0 = pp_5_59_0;
  assign pp_6_59_1 = pp_5_59_1;
  assign pp_6_60_0 = pp_5_60_0;
  assign pp_6_60_1 = pp_5_60_1;
  assign pp_6_61_0 = pp_5_61_0;
  assign pp_6_61_1 = pp_5_61_1;
  assign pp_6_62_0 = pp_5_62_0;
  assign pp_6_62_1 = pp_5_62_1;
  assign pp_7_0_0 = pp_6_0_0;
  assign pp_7_1_0 = pp_6_1_0;
  assign pp_7_1_1 = pp_6_1_1;
  assign pp_7_2_0 = pp_6_2_0;
  assign pp_7_2_1 = pp_6_2_1;
  assign pp_7_3_0 = pp_6_3_0;
  assign pp_7_3_1 = pp_6_3_1;
  assign pp_7_4_0 = pp_6_4_0;
  assign pp_7_4_1 = pp_6_4_1;
  assign pp_7_5_0 = pp_6_5_0;
  assign pp_7_5_1 = pp_6_5_1;
  assign pp_7_6_0 = pp_6_6_0;
  assign pp_7_6_1 = pp_6_6_1;
  assign pp_7_6_2 = pp_6_6_2;
  assign pp_7_7_0 = pp_6_7_0;
  assign pp_7_8_0 = pp_6_8_0;
  assign pp_7_8_1 = pp_6_8_1;
  assign pp_7_9_0 = pp_6_9_0;
  assign pp_7_9_1 = pp_6_9_1;
  assign pp_7_10_0 = pp_6_10_0;
  assign pp_7_10_1 = pp_6_10_1;
  MG_FA fa_6_11_0(
    .a(pp_6_11_0),
    .b(pp_6_11_1),
    .cin(pp_6_11_2),
    .sum(pp_7_11_0),
    .cout(pp_7_12_0)
  );

  assign pp_7_11_1 = pp_6_11_3;
  assign pp_7_12_1 = pp_6_12_0;
  assign pp_7_13_0 = pp_6_13_0;
  assign pp_7_13_1 = pp_6_13_1;
  MG_HA ha_6_14_0(
    .a(pp_6_14_0),
    .b(pp_6_14_1),
    .sum(pp_7_14_0),
    .cout(pp_7_15_0)
  );

  assign pp_7_14_1 = pp_6_14_2;
  assign pp_7_15_1 = pp_6_15_0;
  MG_HA ha_6_16_0(
    .a(pp_6_16_0),
    .b(pp_6_16_1),
    .sum(pp_7_16_0),
    .cout(pp_7_17_0)
  );

  assign pp_7_16_1 = pp_6_16_2;
  assign pp_7_17_1 = pp_6_17_0;
  assign pp_7_17_2 = pp_6_17_1;
  assign pp_7_17_3 = pp_6_17_2;
  assign pp_7_18_0 = pp_6_18_0;
  assign pp_7_18_1 = pp_6_18_1;
  MG_FA fa_6_19_0(
    .a(pp_6_19_0),
    .b(pp_6_19_1),
    .cin(pp_6_19_2),
    .sum(pp_7_19_0),
    .cout(pp_7_20_0)
  );

  assign pp_7_20_1 = pp_6_20_0;
  assign pp_7_20_2 = pp_6_20_1;
  assign pp_7_20_3 = pp_6_20_2;
  assign pp_7_21_0 = pp_6_21_0;
  assign pp_7_21_1 = pp_6_21_1;
  assign pp_7_21_2 = pp_6_21_2;
  MG_HA ha_6_22_0(
    .a(pp_6_22_0),
    .b(pp_6_22_1),
    .sum(pp_7_22_0),
    .cout(pp_7_23_0)
  );

  MG_FA fa_6_23_0(
    .a(pp_6_23_0),
    .b(pp_6_23_1),
    .cin(pp_6_23_2),
    .sum(pp_7_23_1),
    .cout(pp_7_24_0)
  );

  assign pp_7_23_2 = pp_6_23_3;
  MG_FA fa_6_24_0(
    .a(pp_6_24_0),
    .b(pp_6_24_1),
    .cin(pp_6_24_2),
    .sum(pp_7_24_1),
    .cout(pp_7_25_0)
  );

  MG_FA fa_6_25_0(
    .a(pp_6_25_0),
    .b(pp_6_25_1),
    .cin(pp_6_25_2),
    .sum(pp_7_25_1),
    .cout(pp_7_26_0)
  );

  assign pp_7_25_2 = pp_6_25_3;
  MG_FA fa_6_26_0(
    .a(pp_6_26_0),
    .b(pp_6_26_1),
    .cin(pp_6_26_2),
    .sum(pp_7_26_1),
    .cout(pp_7_27_0)
  );

  assign pp_7_26_2 = pp_6_26_3;
  MG_FA fa_6_27_0(
    .a(pp_6_27_0),
    .b(pp_6_27_1),
    .cin(pp_6_27_2),
    .sum(pp_7_27_1),
    .cout(pp_7_28_0)
  );

  MG_HA ha_6_27_1(
    .a(pp_6_27_3),
    .b(pp_6_27_4),
    .sum(pp_7_27_2),
    .cout(pp_7_28_1)
  );

  MG_HA ha_6_28_0(
    .a(pp_6_28_0),
    .b(pp_6_28_1),
    .sum(pp_7_28_2),
    .cout(pp_7_29_0)
  );

  MG_FA fa_6_29_0(
    .a(pp_6_29_0),
    .b(pp_6_29_1),
    .cin(pp_6_29_2),
    .sum(pp_7_29_1),
    .cout(pp_7_30_0)
  );

  assign pp_7_29_2 = pp_6_29_3;
  MG_HA ha_6_30_0(
    .a(pp_6_30_0),
    .b(pp_6_30_1),
    .sum(pp_7_30_1),
    .cout(pp_7_31_0)
  );

  assign pp_7_30_2 = pp_6_30_2;
  MG_HA ha_6_31_0(
    .a(pp_6_31_0),
    .b(pp_6_31_1),
    .sum(pp_7_31_1),
    .cout(pp_7_32_0)
  );

  assign pp_7_31_2 = pp_6_31_2;
  MG_FA fa_6_32_0(
    .a(pp_6_32_0),
    .b(pp_6_32_1),
    .cin(pp_6_32_2),
    .sum(pp_7_32_1),
    .cout(pp_7_33_0)
  );

  MG_HA ha_6_32_1(
    .a(pp_6_32_3),
    .b(pp_6_32_4),
    .sum(pp_7_32_2),
    .cout(pp_7_33_1)
  );

  MG_FA fa_6_33_0(
    .a(pp_6_33_0),
    .b(pp_6_33_1),
    .cin(pp_6_33_2),
    .sum(pp_7_33_2),
    .cout(pp_7_34_0)
  );

  MG_FA fa_6_34_0(
    .a(pp_6_34_0),
    .b(pp_6_34_1),
    .cin(pp_6_34_2),
    .sum(pp_7_34_1),
    .cout(pp_7_35_0)
  );

  assign pp_7_34_2 = pp_6_34_3;
  MG_FA fa_6_35_0(
    .a(pp_6_35_0),
    .b(pp_6_35_1),
    .cin(pp_6_35_2),
    .sum(pp_7_35_1),
    .cout(pp_7_36_0)
  );

  assign pp_7_35_2 = pp_6_35_3;
  MG_FA fa_6_36_0(
    .a(pp_6_36_0),
    .b(pp_6_36_1),
    .cin(pp_6_36_2),
    .sum(pp_7_36_1),
    .cout(pp_7_37_0)
  );

  assign pp_7_36_2 = pp_6_36_3;
  MG_FA fa_6_37_0(
    .a(pp_6_37_0),
    .b(pp_6_37_1),
    .cin(pp_6_37_2),
    .sum(pp_7_37_1),
    .cout(pp_7_38_0)
  );

  assign pp_7_37_2 = pp_6_37_3;
  MG_FA fa_6_38_0(
    .a(pp_6_38_0),
    .b(pp_6_38_1),
    .cin(pp_6_38_2),
    .sum(pp_7_38_1),
    .cout(pp_7_39_0)
  );

  assign pp_7_38_2 = pp_6_38_3;
  MG_FA fa_6_39_0(
    .a(pp_6_39_0),
    .b(pp_6_39_1),
    .cin(pp_6_39_2),
    .sum(pp_7_39_1),
    .cout(pp_7_40_0)
  );

  assign pp_7_39_2 = pp_6_39_3;
  assign pp_7_40_1 = pp_6_40_0;
  assign pp_7_40_2 = pp_6_40_1;
  MG_FA fa_6_41_0(
    .a(pp_6_41_0),
    .b(pp_6_41_1),
    .cin(pp_6_41_2),
    .sum(pp_7_41_0),
    .cout(pp_7_42_0)
  );

  MG_FA fa_6_41_1(
    .a(pp_6_41_3),
    .b(pp_6_41_4),
    .cin(pp_6_41_5),
    .sum(pp_7_41_1),
    .cout(pp_7_42_1)
  );

  assign pp_7_41_2 = pp_6_41_6;
  MG_FA fa_6_42_0(
    .a(pp_6_42_0),
    .b(pp_6_42_1),
    .cin(pp_6_42_2),
    .sum(pp_7_42_2),
    .cout(pp_7_43_0)
  );

  assign pp_7_43_1 = pp_6_43_0;
  assign pp_7_43_2 = pp_6_43_1;
  MG_FA fa_6_44_0(
    .a(pp_6_44_0),
    .b(pp_6_44_1),
    .cin(pp_6_44_2),
    .sum(pp_7_44_0),
    .cout(pp_7_45_0)
  );

  MG_FA fa_6_45_0(
    .a(pp_6_45_0),
    .b(pp_6_45_1),
    .cin(pp_6_45_2),
    .sum(pp_7_45_1),
    .cout(pp_7_46_0)
  );

  assign pp_7_45_2 = pp_6_45_3;
  assign pp_7_45_3 = pp_6_45_4;
  assign pp_7_46_1 = pp_6_46_0;
  assign pp_7_46_2 = pp_6_46_1;
  MG_FA fa_6_47_0(
    .a(pp_6_47_0),
    .b(pp_6_47_1),
    .cin(pp_6_47_2),
    .sum(pp_7_47_0),
    .cout(pp_7_48_0)
  );

  MG_FA fa_6_48_0(
    .a(pp_6_48_0),
    .b(pp_6_48_1),
    .cin(pp_6_48_2),
    .sum(pp_7_48_1),
    .cout(pp_7_49_0)
  );

  assign pp_7_49_1 = pp_6_49_0;
  assign pp_7_49_2 = pp_6_49_1;
  assign pp_7_49_3 = pp_6_49_2;
  assign pp_7_50_0 = pp_6_50_0;
  assign pp_7_50_1 = pp_6_50_1;
  assign pp_7_50_2 = pp_6_50_2;
  MG_FA fa_6_51_0(
    .a(pp_6_51_0),
    .b(pp_6_51_1),
    .cin(pp_6_51_2),
    .sum(pp_7_51_0),
    .cout(pp_7_52_0)
  );

  MG_FA fa_6_52_0(
    .a(pp_6_52_0),
    .b(pp_6_52_1),
    .cin(pp_6_52_2),
    .sum(pp_7_52_1),
    .cout(pp_7_53_0)
  );

  assign pp_7_53_1 = pp_6_53_0;
  assign pp_7_53_2 = pp_6_53_1;
  assign pp_7_53_3 = pp_6_53_2;
  assign pp_7_54_0 = pp_6_54_0;
  assign pp_7_55_0 = pp_6_55_0;
  assign pp_7_55_1 = pp_6_55_1;
  assign pp_7_56_0 = pp_6_56_0;
  assign pp_7_56_1 = pp_6_56_1;
  assign pp_7_57_0 = pp_6_57_0;
  assign pp_7_57_1 = pp_6_57_1;
  assign pp_7_58_0 = pp_6_58_0;
  assign pp_7_58_1 = pp_6_58_1;
  assign pp_7_59_0 = pp_6_59_0;
  assign pp_7_59_1 = pp_6_59_1;
  assign pp_7_60_0 = pp_6_60_0;
  assign pp_7_60_1 = pp_6_60_1;
  assign pp_7_61_0 = pp_6_61_0;
  assign pp_7_61_1 = pp_6_61_1;
  assign pp_7_62_0 = pp_6_62_0;
  assign pp_7_62_1 = pp_6_62_1;
  assign pp_8_0_0 = pp_7_0_0;
  assign pp_8_1_0 = pp_7_1_0;
  assign pp_8_1_1 = pp_7_1_1;
  assign pp_8_2_0 = pp_7_2_0;
  assign pp_8_2_1 = pp_7_2_1;
  assign pp_8_3_0 = pp_7_3_0;
  assign pp_8_3_1 = pp_7_3_1;
  assign pp_8_4_0 = pp_7_4_0;
  assign pp_8_4_1 = pp_7_4_1;
  assign pp_8_5_0 = pp_7_5_0;
  assign pp_8_5_1 = pp_7_5_1;
  MG_HA ha_7_6_0(
    .a(pp_7_6_0),
    .b(pp_7_6_1),
    .sum(pp_8_6_0),
    .cout(pp_8_7_0)
  );

  assign pp_8_6_1 = pp_7_6_2;
  assign pp_8_7_1 = pp_7_7_0;
  assign pp_8_8_0 = pp_7_8_0;
  assign pp_8_8_1 = pp_7_8_1;
  assign pp_8_9_0 = pp_7_9_0;
  assign pp_8_9_1 = pp_7_9_1;
  assign pp_8_10_0 = pp_7_10_0;
  assign pp_8_10_1 = pp_7_10_1;
  assign pp_8_11_0 = pp_7_11_0;
  assign pp_8_11_1 = pp_7_11_1;
  assign pp_8_12_0 = pp_7_12_0;
  assign pp_8_12_1 = pp_7_12_1;
  assign pp_8_13_0 = pp_7_13_0;
  assign pp_8_13_1 = pp_7_13_1;
  assign pp_8_14_0 = pp_7_14_0;
  assign pp_8_14_1 = pp_7_14_1;
  assign pp_8_15_0 = pp_7_15_0;
  assign pp_8_15_1 = pp_7_15_1;
  assign pp_8_16_0 = pp_7_16_0;
  assign pp_8_16_1 = pp_7_16_1;
  MG_FA fa_7_17_0(
    .a(pp_7_17_0),
    .b(pp_7_17_1),
    .cin(pp_7_17_2),
    .sum(pp_8_17_0),
    .cout(pp_8_18_0)
  );

  assign pp_8_17_1 = pp_7_17_3;
  MG_HA ha_7_18_0(
    .a(pp_7_18_0),
    .b(pp_7_18_1),
    .sum(pp_8_18_1),
    .cout(pp_8_19_0)
  );

  assign pp_8_19_1 = pp_7_19_0;
  MG_FA fa_7_20_0(
    .a(pp_7_20_0),
    .b(pp_7_20_1),
    .cin(pp_7_20_2),
    .sum(pp_8_20_0),
    .cout(pp_8_21_0)
  );

  assign pp_8_20_1 = pp_7_20_3;
  MG_FA fa_7_21_0(
    .a(pp_7_21_0),
    .b(pp_7_21_1),
    .cin(pp_7_21_2),
    .sum(pp_8_21_1),
    .cout(pp_8_22_0)
  );

  assign pp_8_22_1 = pp_7_22_0;
  MG_HA ha_7_23_0(
    .a(pp_7_23_0),
    .b(pp_7_23_1),
    .sum(pp_8_23_0),
    .cout(pp_8_24_0)
  );

  assign pp_8_23_1 = pp_7_23_2;
  MG_HA ha_7_24_0(
    .a(pp_7_24_0),
    .b(pp_7_24_1),
    .sum(pp_8_24_1),
    .cout(pp_8_25_0)
  );

  MG_FA fa_7_25_0(
    .a(pp_7_25_0),
    .b(pp_7_25_1),
    .cin(pp_7_25_2),
    .sum(pp_8_25_1),
    .cout(pp_8_26_0)
  );

  MG_FA fa_7_26_0(
    .a(pp_7_26_0),
    .b(pp_7_26_1),
    .cin(pp_7_26_2),
    .sum(pp_8_26_1),
    .cout(pp_8_27_0)
  );

  MG_FA fa_7_27_0(
    .a(pp_7_27_0),
    .b(pp_7_27_1),
    .cin(pp_7_27_2),
    .sum(pp_8_27_1),
    .cout(pp_8_28_0)
  );

  MG_FA fa_7_28_0(
    .a(pp_7_28_0),
    .b(pp_7_28_1),
    .cin(pp_7_28_2),
    .sum(pp_8_28_1),
    .cout(pp_8_29_0)
  );

  MG_FA fa_7_29_0(
    .a(pp_7_29_0),
    .b(pp_7_29_1),
    .cin(pp_7_29_2),
    .sum(pp_8_29_1),
    .cout(pp_8_30_0)
  );

  MG_FA fa_7_30_0(
    .a(pp_7_30_0),
    .b(pp_7_30_1),
    .cin(pp_7_30_2),
    .sum(pp_8_30_1),
    .cout(pp_8_31_0)
  );

  MG_FA fa_7_31_0(
    .a(pp_7_31_0),
    .b(pp_7_31_1),
    .cin(pp_7_31_2),
    .sum(pp_8_31_1),
    .cout(pp_8_32_0)
  );

  MG_FA fa_7_32_0(
    .a(pp_7_32_0),
    .b(pp_7_32_1),
    .cin(pp_7_32_2),
    .sum(pp_8_32_1),
    .cout(pp_8_33_0)
  );

  MG_FA fa_7_33_0(
    .a(pp_7_33_0),
    .b(pp_7_33_1),
    .cin(pp_7_33_2),
    .sum(pp_8_33_1),
    .cout(pp_8_34_0)
  );

  MG_FA fa_7_34_0(
    .a(pp_7_34_0),
    .b(pp_7_34_1),
    .cin(pp_7_34_2),
    .sum(pp_8_34_1),
    .cout(pp_8_35_0)
  );

  MG_FA fa_7_35_0(
    .a(pp_7_35_0),
    .b(pp_7_35_1),
    .cin(pp_7_35_2),
    .sum(pp_8_35_1),
    .cout(pp_8_36_0)
  );

  MG_FA fa_7_36_0(
    .a(pp_7_36_0),
    .b(pp_7_36_1),
    .cin(pp_7_36_2),
    .sum(pp_8_36_1),
    .cout(pp_8_37_0)
  );

  MG_FA fa_7_37_0(
    .a(pp_7_37_0),
    .b(pp_7_37_1),
    .cin(pp_7_37_2),
    .sum(pp_8_37_1),
    .cout(pp_8_38_0)
  );

  MG_FA fa_7_38_0(
    .a(pp_7_38_0),
    .b(pp_7_38_1),
    .cin(pp_7_38_2),
    .sum(pp_8_38_1),
    .cout(pp_8_39_0)
  );

  MG_FA fa_7_39_0(
    .a(pp_7_39_0),
    .b(pp_7_39_1),
    .cin(pp_7_39_2),
    .sum(pp_8_39_1),
    .cout(pp_8_40_0)
  );

  MG_FA fa_7_40_0(
    .a(pp_7_40_0),
    .b(pp_7_40_1),
    .cin(pp_7_40_2),
    .sum(pp_8_40_1),
    .cout(pp_8_41_0)
  );

  MG_FA fa_7_41_0(
    .a(pp_7_41_0),
    .b(pp_7_41_1),
    .cin(pp_7_41_2),
    .sum(pp_8_41_1),
    .cout(pp_8_42_0)
  );

  MG_FA fa_7_42_0(
    .a(pp_7_42_0),
    .b(pp_7_42_1),
    .cin(pp_7_42_2),
    .sum(pp_8_42_1),
    .cout(pp_8_43_0)
  );

  MG_FA fa_7_43_0(
    .a(pp_7_43_0),
    .b(pp_7_43_1),
    .cin(pp_7_43_2),
    .sum(pp_8_43_1),
    .cout(pp_8_44_0)
  );

  assign pp_8_44_1 = pp_7_44_0;
  MG_FA fa_7_45_0(
    .a(pp_7_45_0),
    .b(pp_7_45_1),
    .cin(pp_7_45_2),
    .sum(pp_8_45_0),
    .cout(pp_8_46_0)
  );

  assign pp_8_45_1 = pp_7_45_3;
  MG_FA fa_7_46_0(
    .a(pp_7_46_0),
    .b(pp_7_46_1),
    .cin(pp_7_46_2),
    .sum(pp_8_46_1),
    .cout(pp_8_47_0)
  );

  assign pp_8_47_1 = pp_7_47_0;
  assign pp_8_48_0 = pp_7_48_0;
  assign pp_8_48_1 = pp_7_48_1;
  MG_FA fa_7_49_0(
    .a(pp_7_49_0),
    .b(pp_7_49_1),
    .cin(pp_7_49_2),
    .sum(pp_8_49_0),
    .cout(pp_8_50_0)
  );

  assign pp_8_49_1 = pp_7_49_3;
  MG_FA fa_7_50_0(
    .a(pp_7_50_0),
    .b(pp_7_50_1),
    .cin(pp_7_50_2),
    .sum(pp_8_50_1),
    .cout(pp_8_51_0)
  );

  assign pp_8_51_1 = pp_7_51_0;
  assign pp_8_52_0 = pp_7_52_0;
  assign pp_8_52_1 = pp_7_52_1;
  MG_FA fa_7_53_0(
    .a(pp_7_53_0),
    .b(pp_7_53_1),
    .cin(pp_7_53_2),
    .sum(pp_8_53_0),
    .cout(pp_8_54_0)
  );

  assign pp_8_53_1 = pp_7_53_3;
  assign pp_8_54_1 = pp_7_54_0;
  assign pp_8_55_0 = pp_7_55_0;
  assign pp_8_55_1 = pp_7_55_1;
  assign pp_8_56_0 = pp_7_56_0;
  assign pp_8_56_1 = pp_7_56_1;
  assign pp_8_57_0 = pp_7_57_0;
  assign pp_8_57_1 = pp_7_57_1;
  assign pp_8_58_0 = pp_7_58_0;
  assign pp_8_58_1 = pp_7_58_1;
  assign pp_8_59_0 = pp_7_59_0;
  assign pp_8_59_1 = pp_7_59_1;
  assign pp_8_60_0 = pp_7_60_0;
  assign pp_8_60_1 = pp_7_60_1;
  assign pp_8_61_0 = pp_7_61_0;
  assign pp_8_61_1 = pp_7_61_1;
  assign pp_8_62_0 = pp_7_62_0;
  assign pp_8_62_1 = pp_7_62_1;
  wire [61:0] cta;
  wire [61:0] ctb;
  wire [61:0] cts;
  wire ctc;

  MG_CPA cpa(
 .a(cta), .b(ctb), .sum(cts), .cout(ctc)
  );

  assign cta[0] = pp_8_1_0;
  assign ctb[0] = pp_8_1_1;
  assign cta[1] = pp_8_2_0;
  assign ctb[1] = pp_8_2_1;
  assign cta[2] = pp_8_3_0;
  assign ctb[2] = pp_8_3_1;
  assign cta[3] = pp_8_4_0;
  assign ctb[3] = pp_8_4_1;
  assign cta[4] = pp_8_5_0;
  assign ctb[4] = pp_8_5_1;
  assign cta[5] = pp_8_6_0;
  assign ctb[5] = pp_8_6_1;
  assign cta[6] = pp_8_7_0;
  assign ctb[6] = pp_8_7_1;
  assign cta[7] = pp_8_8_0;
  assign ctb[7] = pp_8_8_1;
  assign cta[8] = pp_8_9_0;
  assign ctb[8] = pp_8_9_1;
  assign cta[9] = pp_8_10_0;
  assign ctb[9] = pp_8_10_1;
  assign cta[10] = pp_8_11_0;
  assign ctb[10] = pp_8_11_1;
  assign cta[11] = pp_8_12_0;
  assign ctb[11] = pp_8_12_1;
  assign cta[12] = pp_8_13_0;
  assign ctb[12] = pp_8_13_1;
  assign cta[13] = pp_8_14_0;
  assign ctb[13] = pp_8_14_1;
  assign cta[14] = pp_8_15_0;
  assign ctb[14] = pp_8_15_1;
  assign cta[15] = pp_8_16_0;
  assign ctb[15] = pp_8_16_1;
  assign cta[16] = pp_8_17_0;
  assign ctb[16] = pp_8_17_1;
  assign cta[17] = pp_8_18_0;
  assign ctb[17] = pp_8_18_1;
  assign cta[18] = pp_8_19_0;
  assign ctb[18] = pp_8_19_1;
  assign cta[19] = pp_8_20_0;
  assign ctb[19] = pp_8_20_1;
  assign cta[20] = pp_8_21_0;
  assign ctb[20] = pp_8_21_1;
  assign cta[21] = pp_8_22_0;
  assign ctb[21] = pp_8_22_1;
  assign cta[22] = pp_8_23_0;
  assign ctb[22] = pp_8_23_1;
  assign cta[23] = pp_8_24_0;
  assign ctb[23] = pp_8_24_1;
  assign cta[24] = pp_8_25_0;
  assign ctb[24] = pp_8_25_1;
  assign cta[25] = pp_8_26_0;
  assign ctb[25] = pp_8_26_1;
  assign cta[26] = pp_8_27_0;
  assign ctb[26] = pp_8_27_1;
  assign cta[27] = pp_8_28_0;
  assign ctb[27] = pp_8_28_1;
  assign cta[28] = pp_8_29_0;
  assign ctb[28] = pp_8_29_1;
  assign cta[29] = pp_8_30_0;
  assign ctb[29] = pp_8_30_1;
  assign cta[30] = pp_8_31_0;
  assign ctb[30] = pp_8_31_1;
  assign cta[31] = pp_8_32_0;
  assign ctb[31] = pp_8_32_1;
  assign cta[32] = pp_8_33_0;
  assign ctb[32] = pp_8_33_1;
  assign cta[33] = pp_8_34_0;
  assign ctb[33] = pp_8_34_1;
  assign cta[34] = pp_8_35_0;
  assign ctb[34] = pp_8_35_1;
  assign cta[35] = pp_8_36_0;
  assign ctb[35] = pp_8_36_1;
  assign cta[36] = pp_8_37_0;
  assign ctb[36] = pp_8_37_1;
  assign cta[37] = pp_8_38_0;
  assign ctb[37] = pp_8_38_1;
  assign cta[38] = pp_8_39_0;
  assign ctb[38] = pp_8_39_1;
  assign cta[39] = pp_8_40_0;
  assign ctb[39] = pp_8_40_1;
  assign cta[40] = pp_8_41_0;
  assign ctb[40] = pp_8_41_1;
  assign cta[41] = pp_8_42_0;
  assign ctb[41] = pp_8_42_1;
  assign cta[42] = pp_8_43_0;
  assign ctb[42] = pp_8_43_1;
  assign cta[43] = pp_8_44_0;
  assign ctb[43] = pp_8_44_1;
  assign cta[44] = pp_8_45_0;
  assign ctb[44] = pp_8_45_1;
  assign cta[45] = pp_8_46_0;
  assign ctb[45] = pp_8_46_1;
  assign cta[46] = pp_8_47_0;
  assign ctb[46] = pp_8_47_1;
  assign cta[47] = pp_8_48_0;
  assign ctb[47] = pp_8_48_1;
  assign cta[48] = pp_8_49_0;
  assign ctb[48] = pp_8_49_1;
  assign cta[49] = pp_8_50_0;
  assign ctb[49] = pp_8_50_1;
  assign cta[50] = pp_8_51_0;
  assign ctb[50] = pp_8_51_1;
  assign cta[51] = pp_8_52_0;
  assign ctb[51] = pp_8_52_1;
  assign cta[52] = pp_8_53_0;
  assign ctb[52] = pp_8_53_1;
  assign cta[53] = pp_8_54_0;
  assign ctb[53] = pp_8_54_1;
  assign cta[54] = pp_8_55_0;
  assign ctb[54] = pp_8_55_1;
  assign cta[55] = pp_8_56_0;
  assign ctb[55] = pp_8_56_1;
  assign cta[56] = pp_8_57_0;
  assign ctb[56] = pp_8_57_1;
  assign cta[57] = pp_8_58_0;
  assign ctb[57] = pp_8_58_1;
  assign cta[58] = pp_8_59_0;
  assign ctb[58] = pp_8_59_1;
  assign cta[59] = pp_8_60_0;
  assign ctb[59] = pp_8_60_1;
  assign cta[60] = pp_8_61_0;
  assign ctb[60] = pp_8_61_1;
  assign cta[61] = pp_8_62_0;
  assign ctb[61] = pp_8_62_1;
  assign product[0] = pp_8_0_0;
  assign product[62:1] = cts;
  assign product[63] = ctc;
endmodule
