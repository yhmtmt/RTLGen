module MG_CPA(
  input [30:0] a,
  input [30:0] b,
  output [30:0] sum,
  output cout
);

  wire p_0_0;
  wire g_0_0;
 assign p_0_0 = a[0] ^ b[0];
 assign g_0_0 = a[0] & b[0];
  wire p_1_1;
  wire g_1_1;
 assign p_1_1 = a[1] ^ b[1];
 assign g_1_1 = a[1] & b[1];
  wire p_1_0;
  wire g_1_0;
  wire p_2_2;
  wire g_2_2;
 assign p_2_2 = a[2] ^ b[2];
 assign g_2_2 = a[2] & b[2];
  wire p_2_0;
  wire g_2_0;
  wire p_2_1;
  wire g_2_1;
  wire p_3_3;
  wire g_3_3;
 assign p_3_3 = a[3] ^ b[3];
 assign g_3_3 = a[3] & b[3];
  wire p_3_0;
  wire g_3_0;
  wire p_3_1;
  wire g_3_1;
  wire p_3_2;
  wire g_3_2;
  wire p_4_4;
  wire g_4_4;
 assign p_4_4 = a[4] ^ b[4];
 assign g_4_4 = a[4] & b[4];
  wire p_4_0;
  wire g_4_0;
  wire p_4_1;
  wire g_4_1;
  wire p_4_2;
  wire g_4_2;
  wire p_4_3;
  wire g_4_3;
  wire p_5_5;
  wire g_5_5;
 assign p_5_5 = a[5] ^ b[5];
 assign g_5_5 = a[5] & b[5];
  wire p_5_0;
  wire g_5_0;
  wire p_5_1;
  wire g_5_1;
  wire p_5_2;
  wire g_5_2;
  wire p_5_3;
  wire g_5_3;
  wire p_5_4;
  wire g_5_4;
  wire p_6_6;
  wire g_6_6;
 assign p_6_6 = a[6] ^ b[6];
 assign g_6_6 = a[6] & b[6];
  wire p_6_0;
  wire g_6_0;
  wire p_6_1;
  wire g_6_1;
  wire p_6_2;
  wire g_6_2;
  wire p_6_3;
  wire g_6_3;
  wire p_6_4;
  wire g_6_4;
  wire p_6_5;
  wire g_6_5;
  wire p_7_7;
  wire g_7_7;
 assign p_7_7 = a[7] ^ b[7];
 assign g_7_7 = a[7] & b[7];
  wire p_7_0;
  wire g_7_0;
  wire p_7_1;
  wire g_7_1;
  wire p_7_2;
  wire g_7_2;
  wire p_7_3;
  wire g_7_3;
  wire p_7_4;
  wire g_7_4;
  wire p_7_5;
  wire g_7_5;
  wire p_7_6;
  wire g_7_6;
  wire p_8_8;
  wire g_8_8;
 assign p_8_8 = a[8] ^ b[8];
 assign g_8_8 = a[8] & b[8];
  wire p_8_0;
  wire g_8_0;
  wire p_8_1;
  wire g_8_1;
  wire p_8_2;
  wire g_8_2;
  wire p_8_3;
  wire g_8_3;
  wire p_8_4;
  wire g_8_4;
  wire p_8_5;
  wire g_8_5;
  wire p_8_6;
  wire g_8_6;
  wire p_8_7;
  wire g_8_7;
  wire p_9_9;
  wire g_9_9;
 assign p_9_9 = a[9] ^ b[9];
 assign g_9_9 = a[9] & b[9];
  wire p_9_0;
  wire g_9_0;
  wire p_9_1;
  wire g_9_1;
  wire p_9_2;
  wire g_9_2;
  wire p_9_3;
  wire g_9_3;
  wire p_9_4;
  wire g_9_4;
  wire p_9_5;
  wire g_9_5;
  wire p_9_6;
  wire g_9_6;
  wire p_9_7;
  wire g_9_7;
  wire p_9_8;
  wire g_9_8;
  wire p_10_10;
  wire g_10_10;
 assign p_10_10 = a[10] ^ b[10];
 assign g_10_10 = a[10] & b[10];
  wire p_10_0;
  wire g_10_0;
  wire p_10_1;
  wire g_10_1;
  wire p_10_2;
  wire g_10_2;
  wire p_10_3;
  wire g_10_3;
  wire p_10_4;
  wire g_10_4;
  wire p_10_5;
  wire g_10_5;
  wire p_10_6;
  wire g_10_6;
  wire p_10_7;
  wire g_10_7;
  wire p_10_8;
  wire g_10_8;
  wire p_10_9;
  wire g_10_9;
  wire p_11_11;
  wire g_11_11;
 assign p_11_11 = a[11] ^ b[11];
 assign g_11_11 = a[11] & b[11];
  wire p_11_0;
  wire g_11_0;
  wire p_11_1;
  wire g_11_1;
  wire p_11_2;
  wire g_11_2;
  wire p_11_3;
  wire g_11_3;
  wire p_11_4;
  wire g_11_4;
  wire p_11_5;
  wire g_11_5;
  wire p_11_6;
  wire g_11_6;
  wire p_11_7;
  wire g_11_7;
  wire p_11_8;
  wire g_11_8;
  wire p_11_9;
  wire g_11_9;
  wire p_11_10;
  wire g_11_10;
  wire p_12_12;
  wire g_12_12;
 assign p_12_12 = a[12] ^ b[12];
 assign g_12_12 = a[12] & b[12];
  wire p_12_0;
  wire g_12_0;
  wire p_12_1;
  wire g_12_1;
  wire p_12_2;
  wire g_12_2;
  wire p_12_3;
  wire g_12_3;
  wire p_12_4;
  wire g_12_4;
  wire p_12_5;
  wire g_12_5;
  wire p_12_6;
  wire g_12_6;
  wire p_12_7;
  wire g_12_7;
  wire p_12_8;
  wire g_12_8;
  wire p_12_9;
  wire g_12_9;
  wire p_12_10;
  wire g_12_10;
  wire p_12_11;
  wire g_12_11;
  wire p_13_13;
  wire g_13_13;
 assign p_13_13 = a[13] ^ b[13];
 assign g_13_13 = a[13] & b[13];
  wire p_13_0;
  wire g_13_0;
  wire p_13_1;
  wire g_13_1;
  wire p_13_2;
  wire g_13_2;
  wire p_13_3;
  wire g_13_3;
  wire p_13_4;
  wire g_13_4;
  wire p_13_5;
  wire g_13_5;
  wire p_13_6;
  wire g_13_6;
  wire p_13_7;
  wire g_13_7;
  wire p_13_8;
  wire g_13_8;
  wire p_13_9;
  wire g_13_9;
  wire p_13_10;
  wire g_13_10;
  wire p_13_11;
  wire g_13_11;
  wire p_13_12;
  wire g_13_12;
  wire p_14_14;
  wire g_14_14;
 assign p_14_14 = a[14] ^ b[14];
 assign g_14_14 = a[14] & b[14];
  wire p_14_0;
  wire g_14_0;
  wire p_14_1;
  wire g_14_1;
  wire p_14_2;
  wire g_14_2;
  wire p_14_3;
  wire g_14_3;
  wire p_14_4;
  wire g_14_4;
  wire p_14_5;
  wire g_14_5;
  wire p_14_6;
  wire g_14_6;
  wire p_14_7;
  wire g_14_7;
  wire p_14_8;
  wire g_14_8;
  wire p_14_9;
  wire g_14_9;
  wire p_14_10;
  wire g_14_10;
  wire p_14_11;
  wire g_14_11;
  wire p_14_12;
  wire g_14_12;
  wire p_14_13;
  wire g_14_13;
  wire p_15_15;
  wire g_15_15;
 assign p_15_15 = a[15] ^ b[15];
 assign g_15_15 = a[15] & b[15];
  wire p_15_0;
  wire g_15_0;
  wire p_15_1;
  wire g_15_1;
  wire p_15_2;
  wire g_15_2;
  wire p_15_3;
  wire g_15_3;
  wire p_15_4;
  wire g_15_4;
  wire p_15_5;
  wire g_15_5;
  wire p_15_6;
  wire g_15_6;
  wire p_15_7;
  wire g_15_7;
  wire p_15_8;
  wire g_15_8;
  wire p_15_9;
  wire g_15_9;
  wire p_15_10;
  wire g_15_10;
  wire p_15_11;
  wire g_15_11;
  wire p_15_12;
  wire g_15_12;
  wire p_15_13;
  wire g_15_13;
  wire p_15_14;
  wire g_15_14;
  wire p_16_16;
  wire g_16_16;
 assign p_16_16 = a[16] ^ b[16];
 assign g_16_16 = a[16] & b[16];
  wire p_16_0;
  wire g_16_0;
  wire p_16_1;
  wire g_16_1;
  wire p_16_2;
  wire g_16_2;
  wire p_16_3;
  wire g_16_3;
  wire p_16_4;
  wire g_16_4;
  wire p_16_5;
  wire g_16_5;
  wire p_16_6;
  wire g_16_6;
  wire p_16_7;
  wire g_16_7;
  wire p_16_8;
  wire g_16_8;
  wire p_16_9;
  wire g_16_9;
  wire p_16_10;
  wire g_16_10;
  wire p_16_11;
  wire g_16_11;
  wire p_16_12;
  wire g_16_12;
  wire p_16_13;
  wire g_16_13;
  wire p_16_14;
  wire g_16_14;
  wire p_16_15;
  wire g_16_15;
  wire p_17_17;
  wire g_17_17;
 assign p_17_17 = a[17] ^ b[17];
 assign g_17_17 = a[17] & b[17];
  wire p_17_0;
  wire g_17_0;
  wire p_17_1;
  wire g_17_1;
  wire p_17_2;
  wire g_17_2;
  wire p_17_3;
  wire g_17_3;
  wire p_17_4;
  wire g_17_4;
  wire p_17_5;
  wire g_17_5;
  wire p_17_6;
  wire g_17_6;
  wire p_17_7;
  wire g_17_7;
  wire p_17_8;
  wire g_17_8;
  wire p_17_9;
  wire g_17_9;
  wire p_17_10;
  wire g_17_10;
  wire p_17_11;
  wire g_17_11;
  wire p_17_12;
  wire g_17_12;
  wire p_17_13;
  wire g_17_13;
  wire p_17_14;
  wire g_17_14;
  wire p_17_15;
  wire g_17_15;
  wire p_17_16;
  wire g_17_16;
  wire p_18_18;
  wire g_18_18;
 assign p_18_18 = a[18] ^ b[18];
 assign g_18_18 = a[18] & b[18];
  wire p_18_0;
  wire g_18_0;
  wire p_18_1;
  wire g_18_1;
  wire p_18_2;
  wire g_18_2;
  wire p_18_3;
  wire g_18_3;
  wire p_18_4;
  wire g_18_4;
  wire p_18_5;
  wire g_18_5;
  wire p_18_6;
  wire g_18_6;
  wire p_18_7;
  wire g_18_7;
  wire p_18_8;
  wire g_18_8;
  wire p_18_9;
  wire g_18_9;
  wire p_18_10;
  wire g_18_10;
  wire p_18_11;
  wire g_18_11;
  wire p_18_12;
  wire g_18_12;
  wire p_18_13;
  wire g_18_13;
  wire p_18_14;
  wire g_18_14;
  wire p_18_15;
  wire g_18_15;
  wire p_18_16;
  wire g_18_16;
  wire p_18_17;
  wire g_18_17;
  wire p_19_19;
  wire g_19_19;
 assign p_19_19 = a[19] ^ b[19];
 assign g_19_19 = a[19] & b[19];
  wire p_19_0;
  wire g_19_0;
  wire p_19_1;
  wire g_19_1;
  wire p_19_2;
  wire g_19_2;
  wire p_19_3;
  wire g_19_3;
  wire p_19_4;
  wire g_19_4;
  wire p_19_5;
  wire g_19_5;
  wire p_19_6;
  wire g_19_6;
  wire p_19_7;
  wire g_19_7;
  wire p_19_8;
  wire g_19_8;
  wire p_19_9;
  wire g_19_9;
  wire p_19_10;
  wire g_19_10;
  wire p_19_11;
  wire g_19_11;
  wire p_19_12;
  wire g_19_12;
  wire p_19_13;
  wire g_19_13;
  wire p_19_14;
  wire g_19_14;
  wire p_19_15;
  wire g_19_15;
  wire p_19_16;
  wire g_19_16;
  wire p_19_17;
  wire g_19_17;
  wire p_19_18;
  wire g_19_18;
  wire p_20_20;
  wire g_20_20;
 assign p_20_20 = a[20] ^ b[20];
 assign g_20_20 = a[20] & b[20];
  wire p_20_0;
  wire g_20_0;
  wire p_20_1;
  wire g_20_1;
  wire p_20_2;
  wire g_20_2;
  wire p_20_3;
  wire g_20_3;
  wire p_20_4;
  wire g_20_4;
  wire p_20_5;
  wire g_20_5;
  wire p_20_6;
  wire g_20_6;
  wire p_20_7;
  wire g_20_7;
  wire p_20_8;
  wire g_20_8;
  wire p_20_9;
  wire g_20_9;
  wire p_20_10;
  wire g_20_10;
  wire p_20_11;
  wire g_20_11;
  wire p_20_12;
  wire g_20_12;
  wire p_20_13;
  wire g_20_13;
  wire p_20_14;
  wire g_20_14;
  wire p_20_15;
  wire g_20_15;
  wire p_20_16;
  wire g_20_16;
  wire p_20_17;
  wire g_20_17;
  wire p_20_18;
  wire g_20_18;
  wire p_20_19;
  wire g_20_19;
  wire p_21_21;
  wire g_21_21;
 assign p_21_21 = a[21] ^ b[21];
 assign g_21_21 = a[21] & b[21];
  wire p_21_0;
  wire g_21_0;
  wire p_21_1;
  wire g_21_1;
  wire p_21_2;
  wire g_21_2;
  wire p_21_3;
  wire g_21_3;
  wire p_21_4;
  wire g_21_4;
  wire p_21_5;
  wire g_21_5;
  wire p_21_6;
  wire g_21_6;
  wire p_21_7;
  wire g_21_7;
  wire p_21_8;
  wire g_21_8;
  wire p_21_9;
  wire g_21_9;
  wire p_21_10;
  wire g_21_10;
  wire p_21_11;
  wire g_21_11;
  wire p_21_12;
  wire g_21_12;
  wire p_21_13;
  wire g_21_13;
  wire p_21_14;
  wire g_21_14;
  wire p_21_15;
  wire g_21_15;
  wire p_21_16;
  wire g_21_16;
  wire p_21_17;
  wire g_21_17;
  wire p_21_18;
  wire g_21_18;
  wire p_21_19;
  wire g_21_19;
  wire p_21_20;
  wire g_21_20;
  wire p_22_22;
  wire g_22_22;
 assign p_22_22 = a[22] ^ b[22];
 assign g_22_22 = a[22] & b[22];
  wire p_22_0;
  wire g_22_0;
  wire p_22_1;
  wire g_22_1;
  wire p_22_2;
  wire g_22_2;
  wire p_22_3;
  wire g_22_3;
  wire p_22_4;
  wire g_22_4;
  wire p_22_5;
  wire g_22_5;
  wire p_22_6;
  wire g_22_6;
  wire p_22_7;
  wire g_22_7;
  wire p_22_8;
  wire g_22_8;
  wire p_22_9;
  wire g_22_9;
  wire p_22_10;
  wire g_22_10;
  wire p_22_11;
  wire g_22_11;
  wire p_22_12;
  wire g_22_12;
  wire p_22_13;
  wire g_22_13;
  wire p_22_14;
  wire g_22_14;
  wire p_22_15;
  wire g_22_15;
  wire p_22_16;
  wire g_22_16;
  wire p_22_17;
  wire g_22_17;
  wire p_22_18;
  wire g_22_18;
  wire p_22_19;
  wire g_22_19;
  wire p_22_20;
  wire g_22_20;
  wire p_22_21;
  wire g_22_21;
  wire p_23_23;
  wire g_23_23;
 assign p_23_23 = a[23] ^ b[23];
 assign g_23_23 = a[23] & b[23];
  wire p_23_0;
  wire g_23_0;
  wire p_23_1;
  wire g_23_1;
  wire p_23_2;
  wire g_23_2;
  wire p_23_3;
  wire g_23_3;
  wire p_23_4;
  wire g_23_4;
  wire p_23_5;
  wire g_23_5;
  wire p_23_6;
  wire g_23_6;
  wire p_23_7;
  wire g_23_7;
  wire p_23_8;
  wire g_23_8;
  wire p_23_9;
  wire g_23_9;
  wire p_23_10;
  wire g_23_10;
  wire p_23_11;
  wire g_23_11;
  wire p_23_12;
  wire g_23_12;
  wire p_23_13;
  wire g_23_13;
  wire p_23_14;
  wire g_23_14;
  wire p_23_15;
  wire g_23_15;
  wire p_23_16;
  wire g_23_16;
  wire p_23_17;
  wire g_23_17;
  wire p_23_18;
  wire g_23_18;
  wire p_23_19;
  wire g_23_19;
  wire p_23_20;
  wire g_23_20;
  wire p_23_21;
  wire g_23_21;
  wire p_23_22;
  wire g_23_22;
  wire p_24_24;
  wire g_24_24;
 assign p_24_24 = a[24] ^ b[24];
 assign g_24_24 = a[24] & b[24];
  wire p_24_0;
  wire g_24_0;
  wire p_24_1;
  wire g_24_1;
  wire p_24_2;
  wire g_24_2;
  wire p_24_3;
  wire g_24_3;
  wire p_24_4;
  wire g_24_4;
  wire p_24_5;
  wire g_24_5;
  wire p_24_6;
  wire g_24_6;
  wire p_24_7;
  wire g_24_7;
  wire p_24_8;
  wire g_24_8;
  wire p_24_9;
  wire g_24_9;
  wire p_24_10;
  wire g_24_10;
  wire p_24_11;
  wire g_24_11;
  wire p_24_12;
  wire g_24_12;
  wire p_24_13;
  wire g_24_13;
  wire p_24_14;
  wire g_24_14;
  wire p_24_15;
  wire g_24_15;
  wire p_24_16;
  wire g_24_16;
  wire p_24_17;
  wire g_24_17;
  wire p_24_18;
  wire g_24_18;
  wire p_24_19;
  wire g_24_19;
  wire p_24_20;
  wire g_24_20;
  wire p_24_21;
  wire g_24_21;
  wire p_24_22;
  wire g_24_22;
  wire p_24_23;
  wire g_24_23;
  wire p_25_25;
  wire g_25_25;
 assign p_25_25 = a[25] ^ b[25];
 assign g_25_25 = a[25] & b[25];
  wire p_25_0;
  wire g_25_0;
  wire p_25_1;
  wire g_25_1;
  wire p_25_2;
  wire g_25_2;
  wire p_25_3;
  wire g_25_3;
  wire p_25_4;
  wire g_25_4;
  wire p_25_5;
  wire g_25_5;
  wire p_25_6;
  wire g_25_6;
  wire p_25_7;
  wire g_25_7;
  wire p_25_8;
  wire g_25_8;
  wire p_25_9;
  wire g_25_9;
  wire p_25_10;
  wire g_25_10;
  wire p_25_11;
  wire g_25_11;
  wire p_25_12;
  wire g_25_12;
  wire p_25_13;
  wire g_25_13;
  wire p_25_14;
  wire g_25_14;
  wire p_25_15;
  wire g_25_15;
  wire p_25_16;
  wire g_25_16;
  wire p_25_17;
  wire g_25_17;
  wire p_25_18;
  wire g_25_18;
  wire p_25_19;
  wire g_25_19;
  wire p_25_20;
  wire g_25_20;
  wire p_25_21;
  wire g_25_21;
  wire p_25_22;
  wire g_25_22;
  wire p_25_23;
  wire g_25_23;
  wire p_25_24;
  wire g_25_24;
  wire p_26_26;
  wire g_26_26;
 assign p_26_26 = a[26] ^ b[26];
 assign g_26_26 = a[26] & b[26];
  wire p_26_0;
  wire g_26_0;
  wire p_26_1;
  wire g_26_1;
  wire p_26_2;
  wire g_26_2;
  wire p_26_3;
  wire g_26_3;
  wire p_26_4;
  wire g_26_4;
  wire p_26_5;
  wire g_26_5;
  wire p_26_6;
  wire g_26_6;
  wire p_26_7;
  wire g_26_7;
  wire p_26_8;
  wire g_26_8;
  wire p_26_9;
  wire g_26_9;
  wire p_26_10;
  wire g_26_10;
  wire p_26_11;
  wire g_26_11;
  wire p_26_12;
  wire g_26_12;
  wire p_26_13;
  wire g_26_13;
  wire p_26_14;
  wire g_26_14;
  wire p_26_15;
  wire g_26_15;
  wire p_26_16;
  wire g_26_16;
  wire p_26_17;
  wire g_26_17;
  wire p_26_18;
  wire g_26_18;
  wire p_26_19;
  wire g_26_19;
  wire p_26_20;
  wire g_26_20;
  wire p_26_21;
  wire g_26_21;
  wire p_26_22;
  wire g_26_22;
  wire p_26_23;
  wire g_26_23;
  wire p_26_24;
  wire g_26_24;
  wire p_26_25;
  wire g_26_25;
  wire p_27_27;
  wire g_27_27;
 assign p_27_27 = a[27] ^ b[27];
 assign g_27_27 = a[27] & b[27];
  wire p_27_0;
  wire g_27_0;
  wire p_27_1;
  wire g_27_1;
  wire p_27_2;
  wire g_27_2;
  wire p_27_3;
  wire g_27_3;
  wire p_27_4;
  wire g_27_4;
  wire p_27_5;
  wire g_27_5;
  wire p_27_6;
  wire g_27_6;
  wire p_27_7;
  wire g_27_7;
  wire p_27_8;
  wire g_27_8;
  wire p_27_9;
  wire g_27_9;
  wire p_27_10;
  wire g_27_10;
  wire p_27_11;
  wire g_27_11;
  wire p_27_12;
  wire g_27_12;
  wire p_27_13;
  wire g_27_13;
  wire p_27_14;
  wire g_27_14;
  wire p_27_15;
  wire g_27_15;
  wire p_27_16;
  wire g_27_16;
  wire p_27_17;
  wire g_27_17;
  wire p_27_18;
  wire g_27_18;
  wire p_27_19;
  wire g_27_19;
  wire p_27_20;
  wire g_27_20;
  wire p_27_21;
  wire g_27_21;
  wire p_27_22;
  wire g_27_22;
  wire p_27_23;
  wire g_27_23;
  wire p_27_24;
  wire g_27_24;
  wire p_27_25;
  wire g_27_25;
  wire p_27_26;
  wire g_27_26;
  wire p_28_28;
  wire g_28_28;
 assign p_28_28 = a[28] ^ b[28];
 assign g_28_28 = a[28] & b[28];
  wire p_28_0;
  wire g_28_0;
  wire p_28_1;
  wire g_28_1;
  wire p_28_2;
  wire g_28_2;
  wire p_28_3;
  wire g_28_3;
  wire p_28_4;
  wire g_28_4;
  wire p_28_5;
  wire g_28_5;
  wire p_28_6;
  wire g_28_6;
  wire p_28_7;
  wire g_28_7;
  wire p_28_8;
  wire g_28_8;
  wire p_28_9;
  wire g_28_9;
  wire p_28_10;
  wire g_28_10;
  wire p_28_11;
  wire g_28_11;
  wire p_28_12;
  wire g_28_12;
  wire p_28_13;
  wire g_28_13;
  wire p_28_14;
  wire g_28_14;
  wire p_28_15;
  wire g_28_15;
  wire p_28_16;
  wire g_28_16;
  wire p_28_17;
  wire g_28_17;
  wire p_28_18;
  wire g_28_18;
  wire p_28_19;
  wire g_28_19;
  wire p_28_20;
  wire g_28_20;
  wire p_28_21;
  wire g_28_21;
  wire p_28_22;
  wire g_28_22;
  wire p_28_23;
  wire g_28_23;
  wire p_28_24;
  wire g_28_24;
  wire p_28_25;
  wire g_28_25;
  wire p_28_26;
  wire g_28_26;
  wire p_28_27;
  wire g_28_27;
  wire p_29_29;
  wire g_29_29;
 assign p_29_29 = a[29] ^ b[29];
 assign g_29_29 = a[29] & b[29];
  wire p_29_0;
  wire g_29_0;
  wire p_29_1;
  wire g_29_1;
  wire p_29_2;
  wire g_29_2;
  wire p_29_3;
  wire g_29_3;
  wire p_29_4;
  wire g_29_4;
  wire p_29_5;
  wire g_29_5;
  wire p_29_6;
  wire g_29_6;
  wire p_29_7;
  wire g_29_7;
  wire p_29_8;
  wire g_29_8;
  wire p_29_9;
  wire g_29_9;
  wire p_29_10;
  wire g_29_10;
  wire p_29_11;
  wire g_29_11;
  wire p_29_12;
  wire g_29_12;
  wire p_29_13;
  wire g_29_13;
  wire p_29_14;
  wire g_29_14;
  wire p_29_15;
  wire g_29_15;
  wire p_29_16;
  wire g_29_16;
  wire p_29_17;
  wire g_29_17;
  wire p_29_18;
  wire g_29_18;
  wire p_29_19;
  wire g_29_19;
  wire p_29_20;
  wire g_29_20;
  wire p_29_21;
  wire g_29_21;
  wire p_29_22;
  wire g_29_22;
  wire p_29_23;
  wire g_29_23;
  wire p_29_24;
  wire g_29_24;
  wire p_29_25;
  wire g_29_25;
  wire p_29_26;
  wire g_29_26;
  wire p_29_27;
  wire g_29_27;
  wire p_29_28;
  wire g_29_28;
  wire p_30_30;
  wire g_30_30;
 assign p_30_30 = a[30] ^ b[30];
 assign g_30_30 = a[30] & b[30];
  wire p_30_0;
  wire g_30_0;
  wire p_30_1;
  wire g_30_1;
  wire p_30_2;
  wire g_30_2;
  wire p_30_3;
  wire g_30_3;
  wire p_30_4;
  wire g_30_4;
  wire p_30_5;
  wire g_30_5;
  wire p_30_6;
  wire g_30_6;
  wire p_30_7;
  wire g_30_7;
  wire p_30_8;
  wire g_30_8;
  wire p_30_9;
  wire g_30_9;
  wire p_30_10;
  wire g_30_10;
  wire p_30_11;
  wire g_30_11;
  wire p_30_12;
  wire g_30_12;
  wire p_30_13;
  wire g_30_13;
  wire p_30_14;
  wire g_30_14;
  wire p_30_15;
  wire g_30_15;
  wire p_30_16;
  wire g_30_16;
  wire p_30_17;
  wire g_30_17;
  wire p_30_18;
  wire g_30_18;
  wire p_30_19;
  wire g_30_19;
  wire p_30_20;
  wire g_30_20;
  wire p_30_21;
  wire g_30_21;
  wire p_30_22;
  wire g_30_22;
  wire p_30_23;
  wire g_30_23;
  wire p_30_24;
  wire g_30_24;
  wire p_30_25;
  wire g_30_25;
  wire p_30_26;
  wire g_30_26;
  wire p_30_27;
  wire g_30_27;
  wire p_30_28;
  wire g_30_28;
  wire p_30_29;
  wire g_30_29;
 assign sum[0] = p_0_0;
 assign p_1_0 = p_1_1 & p_0_0;
 assign g_1_0 = g_1_1 | (p_1_1 & g_0_0);
 assign sum[1] = p_1_1^ g_0_0;
 assign p_2_0 = p_2_1 & p_0_0;
 assign g_2_0 = g_2_1 | (p_2_1 & g_0_0);
 assign p_2_1 = p_2_2 & p_1_1;
 assign g_2_1 = g_2_2 | (p_2_2 & g_1_1);
 assign sum[2] = p_2_2^ g_1_0;
 assign p_3_0 = p_3_2 & p_1_0;
 assign g_3_0 = g_3_2 | (p_3_2 & g_1_0);
 assign p_3_1 = p_3_2 & p_1_1;
 assign g_3_1 = g_3_2 | (p_3_2 & g_1_1);
 assign p_3_2 = p_3_3 & p_2_2;
 assign g_3_2 = g_3_3 | (p_3_3 & g_2_2);
 assign sum[3] = p_3_3^ g_2_0;
 assign p_4_0 = p_4_1 & p_0_0;
 assign g_4_0 = g_4_1 | (p_4_1 & g_0_0);
 assign p_4_1 = p_4_3 & p_2_1;
 assign g_4_1 = g_4_3 | (p_4_3 & g_2_1);
 assign p_4_2 = p_4_3 & p_2_2;
 assign g_4_2 = g_4_3 | (p_4_3 & g_2_2);
 assign p_4_3 = p_4_4 & p_3_3;
 assign g_4_3 = g_4_4 | (p_4_4 & g_3_3);
 assign sum[4] = p_4_4^ g_3_0;
 assign p_5_0 = p_5_2 & p_1_0;
 assign g_5_0 = g_5_2 | (p_5_2 & g_1_0);
 assign p_5_1 = p_5_2 & p_1_1;
 assign g_5_1 = g_5_2 | (p_5_2 & g_1_1);
 assign p_5_2 = p_5_4 & p_3_2;
 assign g_5_2 = g_5_4 | (p_5_4 & g_3_2);
 assign p_5_3 = p_5_4 & p_3_3;
 assign g_5_3 = g_5_4 | (p_5_4 & g_3_3);
 assign p_5_4 = p_5_5 & p_4_4;
 assign g_5_4 = g_5_5 | (p_5_5 & g_4_4);
 assign sum[5] = p_5_5^ g_4_0;
 assign p_6_0 = p_6_3 & p_2_0;
 assign g_6_0 = g_6_3 | (p_6_3 & g_2_0);
 assign p_6_1 = p_6_3 & p_2_1;
 assign g_6_1 = g_6_3 | (p_6_3 & g_2_1);
 assign p_6_2 = p_6_3 & p_2_2;
 assign g_6_2 = g_6_3 | (p_6_3 & g_2_2);
 assign p_6_3 = p_6_5 & p_4_3;
 assign g_6_3 = g_6_5 | (p_6_5 & g_4_3);
 assign p_6_4 = p_6_5 & p_4_4;
 assign g_6_4 = g_6_5 | (p_6_5 & g_4_4);
 assign p_6_5 = p_6_6 & p_5_5;
 assign g_6_5 = g_6_6 | (p_6_6 & g_5_5);
 assign sum[6] = p_6_6^ g_5_0;
 assign p_7_0 = p_7_4 & p_3_0;
 assign g_7_0 = g_7_4 | (p_7_4 & g_3_0);
 assign p_7_1 = p_7_4 & p_3_1;
 assign g_7_1 = g_7_4 | (p_7_4 & g_3_1);
 assign p_7_2 = p_7_4 & p_3_2;
 assign g_7_2 = g_7_4 | (p_7_4 & g_3_2);
 assign p_7_3 = p_7_4 & p_3_3;
 assign g_7_3 = g_7_4 | (p_7_4 & g_3_3);
 assign p_7_4 = p_7_6 & p_5_4;
 assign g_7_4 = g_7_6 | (p_7_6 & g_5_4);
 assign p_7_5 = p_7_6 & p_5_5;
 assign g_7_5 = g_7_6 | (p_7_6 & g_5_5);
 assign p_7_6 = p_7_7 & p_6_6;
 assign g_7_6 = g_7_7 | (p_7_7 & g_6_6);
 assign sum[7] = p_7_7^ g_6_0;
 assign p_8_0 = p_8_1 & p_0_0;
 assign g_8_0 = g_8_1 | (p_8_1 & g_0_0);
 assign p_8_1 = p_8_5 & p_4_1;
 assign g_8_1 = g_8_5 | (p_8_5 & g_4_1);
 assign p_8_2 = p_8_5 & p_4_2;
 assign g_8_2 = g_8_5 | (p_8_5 & g_4_2);
 assign p_8_3 = p_8_5 & p_4_3;
 assign g_8_3 = g_8_5 | (p_8_5 & g_4_3);
 assign p_8_4 = p_8_5 & p_4_4;
 assign g_8_4 = g_8_5 | (p_8_5 & g_4_4);
 assign p_8_5 = p_8_7 & p_6_5;
 assign g_8_5 = g_8_7 | (p_8_7 & g_6_5);
 assign p_8_6 = p_8_7 & p_6_6;
 assign g_8_6 = g_8_7 | (p_8_7 & g_6_6);
 assign p_8_7 = p_8_8 & p_7_7;
 assign g_8_7 = g_8_8 | (p_8_8 & g_7_7);
 assign sum[8] = p_8_8^ g_7_0;
 assign p_9_0 = p_9_2 & p_1_0;
 assign g_9_0 = g_9_2 | (p_9_2 & g_1_0);
 assign p_9_1 = p_9_2 & p_1_1;
 assign g_9_1 = g_9_2 | (p_9_2 & g_1_1);
 assign p_9_2 = p_9_6 & p_5_2;
 assign g_9_2 = g_9_6 | (p_9_6 & g_5_2);
 assign p_9_3 = p_9_6 & p_5_3;
 assign g_9_3 = g_9_6 | (p_9_6 & g_5_3);
 assign p_9_4 = p_9_6 & p_5_4;
 assign g_9_4 = g_9_6 | (p_9_6 & g_5_4);
 assign p_9_5 = p_9_6 & p_5_5;
 assign g_9_5 = g_9_6 | (p_9_6 & g_5_5);
 assign p_9_6 = p_9_8 & p_7_6;
 assign g_9_6 = g_9_8 | (p_9_8 & g_7_6);
 assign p_9_7 = p_9_8 & p_7_7;
 assign g_9_7 = g_9_8 | (p_9_8 & g_7_7);
 assign p_9_8 = p_9_9 & p_8_8;
 assign g_9_8 = g_9_9 | (p_9_9 & g_8_8);
 assign sum[9] = p_9_9^ g_8_0;
 assign p_10_0 = p_10_3 & p_2_0;
 assign g_10_0 = g_10_3 | (p_10_3 & g_2_0);
 assign p_10_1 = p_10_3 & p_2_1;
 assign g_10_1 = g_10_3 | (p_10_3 & g_2_1);
 assign p_10_2 = p_10_3 & p_2_2;
 assign g_10_2 = g_10_3 | (p_10_3 & g_2_2);
 assign p_10_3 = p_10_7 & p_6_3;
 assign g_10_3 = g_10_7 | (p_10_7 & g_6_3);
 assign p_10_4 = p_10_7 & p_6_4;
 assign g_10_4 = g_10_7 | (p_10_7 & g_6_4);
 assign p_10_5 = p_10_7 & p_6_5;
 assign g_10_5 = g_10_7 | (p_10_7 & g_6_5);
 assign p_10_6 = p_10_7 & p_6_6;
 assign g_10_6 = g_10_7 | (p_10_7 & g_6_6);
 assign p_10_7 = p_10_9 & p_8_7;
 assign g_10_7 = g_10_9 | (p_10_9 & g_8_7);
 assign p_10_8 = p_10_9 & p_8_8;
 assign g_10_8 = g_10_9 | (p_10_9 & g_8_8);
 assign p_10_9 = p_10_10 & p_9_9;
 assign g_10_9 = g_10_10 | (p_10_10 & g_9_9);
 assign sum[10] = p_10_10^ g_9_0;
 assign p_11_0 = p_11_4 & p_3_0;
 assign g_11_0 = g_11_4 | (p_11_4 & g_3_0);
 assign p_11_1 = p_11_4 & p_3_1;
 assign g_11_1 = g_11_4 | (p_11_4 & g_3_1);
 assign p_11_2 = p_11_4 & p_3_2;
 assign g_11_2 = g_11_4 | (p_11_4 & g_3_2);
 assign p_11_3 = p_11_4 & p_3_3;
 assign g_11_3 = g_11_4 | (p_11_4 & g_3_3);
 assign p_11_4 = p_11_8 & p_7_4;
 assign g_11_4 = g_11_8 | (p_11_8 & g_7_4);
 assign p_11_5 = p_11_8 & p_7_5;
 assign g_11_5 = g_11_8 | (p_11_8 & g_7_5);
 assign p_11_6 = p_11_8 & p_7_6;
 assign g_11_6 = g_11_8 | (p_11_8 & g_7_6);
 assign p_11_7 = p_11_8 & p_7_7;
 assign g_11_7 = g_11_8 | (p_11_8 & g_7_7);
 assign p_11_8 = p_11_10 & p_9_8;
 assign g_11_8 = g_11_10 | (p_11_10 & g_9_8);
 assign p_11_9 = p_11_10 & p_9_9;
 assign g_11_9 = g_11_10 | (p_11_10 & g_9_9);
 assign p_11_10 = p_11_11 & p_10_10;
 assign g_11_10 = g_11_11 | (p_11_11 & g_10_10);
 assign sum[11] = p_11_11^ g_10_0;
 assign p_12_0 = p_12_5 & p_4_0;
 assign g_12_0 = g_12_5 | (p_12_5 & g_4_0);
 assign p_12_1 = p_12_5 & p_4_1;
 assign g_12_1 = g_12_5 | (p_12_5 & g_4_1);
 assign p_12_2 = p_12_5 & p_4_2;
 assign g_12_2 = g_12_5 | (p_12_5 & g_4_2);
 assign p_12_3 = p_12_5 & p_4_3;
 assign g_12_3 = g_12_5 | (p_12_5 & g_4_3);
 assign p_12_4 = p_12_5 & p_4_4;
 assign g_12_4 = g_12_5 | (p_12_5 & g_4_4);
 assign p_12_5 = p_12_9 & p_8_5;
 assign g_12_5 = g_12_9 | (p_12_9 & g_8_5);
 assign p_12_6 = p_12_9 & p_8_6;
 assign g_12_6 = g_12_9 | (p_12_9 & g_8_6);
 assign p_12_7 = p_12_9 & p_8_7;
 assign g_12_7 = g_12_9 | (p_12_9 & g_8_7);
 assign p_12_8 = p_12_9 & p_8_8;
 assign g_12_8 = g_12_9 | (p_12_9 & g_8_8);
 assign p_12_9 = p_12_11 & p_10_9;
 assign g_12_9 = g_12_11 | (p_12_11 & g_10_9);
 assign p_12_10 = p_12_11 & p_10_10;
 assign g_12_10 = g_12_11 | (p_12_11 & g_10_10);
 assign p_12_11 = p_12_12 & p_11_11;
 assign g_12_11 = g_12_12 | (p_12_12 & g_11_11);
 assign sum[12] = p_12_12^ g_11_0;
 assign p_13_0 = p_13_6 & p_5_0;
 assign g_13_0 = g_13_6 | (p_13_6 & g_5_0);
 assign p_13_1 = p_13_6 & p_5_1;
 assign g_13_1 = g_13_6 | (p_13_6 & g_5_1);
 assign p_13_2 = p_13_6 & p_5_2;
 assign g_13_2 = g_13_6 | (p_13_6 & g_5_2);
 assign p_13_3 = p_13_6 & p_5_3;
 assign g_13_3 = g_13_6 | (p_13_6 & g_5_3);
 assign p_13_4 = p_13_6 & p_5_4;
 assign g_13_4 = g_13_6 | (p_13_6 & g_5_4);
 assign p_13_5 = p_13_6 & p_5_5;
 assign g_13_5 = g_13_6 | (p_13_6 & g_5_5);
 assign p_13_6 = p_13_10 & p_9_6;
 assign g_13_6 = g_13_10 | (p_13_10 & g_9_6);
 assign p_13_7 = p_13_10 & p_9_7;
 assign g_13_7 = g_13_10 | (p_13_10 & g_9_7);
 assign p_13_8 = p_13_10 & p_9_8;
 assign g_13_8 = g_13_10 | (p_13_10 & g_9_8);
 assign p_13_9 = p_13_10 & p_9_9;
 assign g_13_9 = g_13_10 | (p_13_10 & g_9_9);
 assign p_13_10 = p_13_12 & p_11_10;
 assign g_13_10 = g_13_12 | (p_13_12 & g_11_10);
 assign p_13_11 = p_13_12 & p_11_11;
 assign g_13_11 = g_13_12 | (p_13_12 & g_11_11);
 assign p_13_12 = p_13_13 & p_12_12;
 assign g_13_12 = g_13_13 | (p_13_13 & g_12_12);
 assign sum[13] = p_13_13^ g_12_0;
 assign p_14_0 = p_14_7 & p_6_0;
 assign g_14_0 = g_14_7 | (p_14_7 & g_6_0);
 assign p_14_1 = p_14_7 & p_6_1;
 assign g_14_1 = g_14_7 | (p_14_7 & g_6_1);
 assign p_14_2 = p_14_7 & p_6_2;
 assign g_14_2 = g_14_7 | (p_14_7 & g_6_2);
 assign p_14_3 = p_14_7 & p_6_3;
 assign g_14_3 = g_14_7 | (p_14_7 & g_6_3);
 assign p_14_4 = p_14_7 & p_6_4;
 assign g_14_4 = g_14_7 | (p_14_7 & g_6_4);
 assign p_14_5 = p_14_7 & p_6_5;
 assign g_14_5 = g_14_7 | (p_14_7 & g_6_5);
 assign p_14_6 = p_14_7 & p_6_6;
 assign g_14_6 = g_14_7 | (p_14_7 & g_6_6);
 assign p_14_7 = p_14_11 & p_10_7;
 assign g_14_7 = g_14_11 | (p_14_11 & g_10_7);
 assign p_14_8 = p_14_11 & p_10_8;
 assign g_14_8 = g_14_11 | (p_14_11 & g_10_8);
 assign p_14_9 = p_14_11 & p_10_9;
 assign g_14_9 = g_14_11 | (p_14_11 & g_10_9);
 assign p_14_10 = p_14_11 & p_10_10;
 assign g_14_10 = g_14_11 | (p_14_11 & g_10_10);
 assign p_14_11 = p_14_13 & p_12_11;
 assign g_14_11 = g_14_13 | (p_14_13 & g_12_11);
 assign p_14_12 = p_14_13 & p_12_12;
 assign g_14_12 = g_14_13 | (p_14_13 & g_12_12);
 assign p_14_13 = p_14_14 & p_13_13;
 assign g_14_13 = g_14_14 | (p_14_14 & g_13_13);
 assign sum[14] = p_14_14^ g_13_0;
 assign p_15_0 = p_15_8 & p_7_0;
 assign g_15_0 = g_15_8 | (p_15_8 & g_7_0);
 assign p_15_1 = p_15_8 & p_7_1;
 assign g_15_1 = g_15_8 | (p_15_8 & g_7_1);
 assign p_15_2 = p_15_8 & p_7_2;
 assign g_15_2 = g_15_8 | (p_15_8 & g_7_2);
 assign p_15_3 = p_15_8 & p_7_3;
 assign g_15_3 = g_15_8 | (p_15_8 & g_7_3);
 assign p_15_4 = p_15_8 & p_7_4;
 assign g_15_4 = g_15_8 | (p_15_8 & g_7_4);
 assign p_15_5 = p_15_8 & p_7_5;
 assign g_15_5 = g_15_8 | (p_15_8 & g_7_5);
 assign p_15_6 = p_15_8 & p_7_6;
 assign g_15_6 = g_15_8 | (p_15_8 & g_7_6);
 assign p_15_7 = p_15_8 & p_7_7;
 assign g_15_7 = g_15_8 | (p_15_8 & g_7_7);
 assign p_15_8 = p_15_12 & p_11_8;
 assign g_15_8 = g_15_12 | (p_15_12 & g_11_8);
 assign p_15_9 = p_15_12 & p_11_9;
 assign g_15_9 = g_15_12 | (p_15_12 & g_11_9);
 assign p_15_10 = p_15_12 & p_11_10;
 assign g_15_10 = g_15_12 | (p_15_12 & g_11_10);
 assign p_15_11 = p_15_12 & p_11_11;
 assign g_15_11 = g_15_12 | (p_15_12 & g_11_11);
 assign p_15_12 = p_15_14 & p_13_12;
 assign g_15_12 = g_15_14 | (p_15_14 & g_13_12);
 assign p_15_13 = p_15_14 & p_13_13;
 assign g_15_13 = g_15_14 | (p_15_14 & g_13_13);
 assign p_15_14 = p_15_15 & p_14_14;
 assign g_15_14 = g_15_15 | (p_15_15 & g_14_14);
 assign sum[15] = p_15_15^ g_14_0;
 assign p_16_0 = p_16_1 & p_0_0;
 assign g_16_0 = g_16_1 | (p_16_1 & g_0_0);
 assign p_16_1 = p_16_9 & p_8_1;
 assign g_16_1 = g_16_9 | (p_16_9 & g_8_1);
 assign p_16_2 = p_16_9 & p_8_2;
 assign g_16_2 = g_16_9 | (p_16_9 & g_8_2);
 assign p_16_3 = p_16_9 & p_8_3;
 assign g_16_3 = g_16_9 | (p_16_9 & g_8_3);
 assign p_16_4 = p_16_9 & p_8_4;
 assign g_16_4 = g_16_9 | (p_16_9 & g_8_4);
 assign p_16_5 = p_16_9 & p_8_5;
 assign g_16_5 = g_16_9 | (p_16_9 & g_8_5);
 assign p_16_6 = p_16_9 & p_8_6;
 assign g_16_6 = g_16_9 | (p_16_9 & g_8_6);
 assign p_16_7 = p_16_9 & p_8_7;
 assign g_16_7 = g_16_9 | (p_16_9 & g_8_7);
 assign p_16_8 = p_16_9 & p_8_8;
 assign g_16_8 = g_16_9 | (p_16_9 & g_8_8);
 assign p_16_9 = p_16_13 & p_12_9;
 assign g_16_9 = g_16_13 | (p_16_13 & g_12_9);
 assign p_16_10 = p_16_13 & p_12_10;
 assign g_16_10 = g_16_13 | (p_16_13 & g_12_10);
 assign p_16_11 = p_16_13 & p_12_11;
 assign g_16_11 = g_16_13 | (p_16_13 & g_12_11);
 assign p_16_12 = p_16_13 & p_12_12;
 assign g_16_12 = g_16_13 | (p_16_13 & g_12_12);
 assign p_16_13 = p_16_15 & p_14_13;
 assign g_16_13 = g_16_15 | (p_16_15 & g_14_13);
 assign p_16_14 = p_16_15 & p_14_14;
 assign g_16_14 = g_16_15 | (p_16_15 & g_14_14);
 assign p_16_15 = p_16_16 & p_15_15;
 assign g_16_15 = g_16_16 | (p_16_16 & g_15_15);
 assign sum[16] = p_16_16^ g_15_0;
 assign p_17_0 = p_17_2 & p_1_0;
 assign g_17_0 = g_17_2 | (p_17_2 & g_1_0);
 assign p_17_1 = p_17_2 & p_1_1;
 assign g_17_1 = g_17_2 | (p_17_2 & g_1_1);
 assign p_17_2 = p_17_10 & p_9_2;
 assign g_17_2 = g_17_10 | (p_17_10 & g_9_2);
 assign p_17_3 = p_17_10 & p_9_3;
 assign g_17_3 = g_17_10 | (p_17_10 & g_9_3);
 assign p_17_4 = p_17_10 & p_9_4;
 assign g_17_4 = g_17_10 | (p_17_10 & g_9_4);
 assign p_17_5 = p_17_10 & p_9_5;
 assign g_17_5 = g_17_10 | (p_17_10 & g_9_5);
 assign p_17_6 = p_17_10 & p_9_6;
 assign g_17_6 = g_17_10 | (p_17_10 & g_9_6);
 assign p_17_7 = p_17_10 & p_9_7;
 assign g_17_7 = g_17_10 | (p_17_10 & g_9_7);
 assign p_17_8 = p_17_10 & p_9_8;
 assign g_17_8 = g_17_10 | (p_17_10 & g_9_8);
 assign p_17_9 = p_17_10 & p_9_9;
 assign g_17_9 = g_17_10 | (p_17_10 & g_9_9);
 assign p_17_10 = p_17_14 & p_13_10;
 assign g_17_10 = g_17_14 | (p_17_14 & g_13_10);
 assign p_17_11 = p_17_14 & p_13_11;
 assign g_17_11 = g_17_14 | (p_17_14 & g_13_11);
 assign p_17_12 = p_17_14 & p_13_12;
 assign g_17_12 = g_17_14 | (p_17_14 & g_13_12);
 assign p_17_13 = p_17_14 & p_13_13;
 assign g_17_13 = g_17_14 | (p_17_14 & g_13_13);
 assign p_17_14 = p_17_16 & p_15_14;
 assign g_17_14 = g_17_16 | (p_17_16 & g_15_14);
 assign p_17_15 = p_17_16 & p_15_15;
 assign g_17_15 = g_17_16 | (p_17_16 & g_15_15);
 assign p_17_16 = p_17_17 & p_16_16;
 assign g_17_16 = g_17_17 | (p_17_17 & g_16_16);
 assign sum[17] = p_17_17^ g_16_0;
 assign p_18_0 = p_18_3 & p_2_0;
 assign g_18_0 = g_18_3 | (p_18_3 & g_2_0);
 assign p_18_1 = p_18_3 & p_2_1;
 assign g_18_1 = g_18_3 | (p_18_3 & g_2_1);
 assign p_18_2 = p_18_3 & p_2_2;
 assign g_18_2 = g_18_3 | (p_18_3 & g_2_2);
 assign p_18_3 = p_18_11 & p_10_3;
 assign g_18_3 = g_18_11 | (p_18_11 & g_10_3);
 assign p_18_4 = p_18_11 & p_10_4;
 assign g_18_4 = g_18_11 | (p_18_11 & g_10_4);
 assign p_18_5 = p_18_11 & p_10_5;
 assign g_18_5 = g_18_11 | (p_18_11 & g_10_5);
 assign p_18_6 = p_18_11 & p_10_6;
 assign g_18_6 = g_18_11 | (p_18_11 & g_10_6);
 assign p_18_7 = p_18_11 & p_10_7;
 assign g_18_7 = g_18_11 | (p_18_11 & g_10_7);
 assign p_18_8 = p_18_11 & p_10_8;
 assign g_18_8 = g_18_11 | (p_18_11 & g_10_8);
 assign p_18_9 = p_18_11 & p_10_9;
 assign g_18_9 = g_18_11 | (p_18_11 & g_10_9);
 assign p_18_10 = p_18_11 & p_10_10;
 assign g_18_10 = g_18_11 | (p_18_11 & g_10_10);
 assign p_18_11 = p_18_15 & p_14_11;
 assign g_18_11 = g_18_15 | (p_18_15 & g_14_11);
 assign p_18_12 = p_18_15 & p_14_12;
 assign g_18_12 = g_18_15 | (p_18_15 & g_14_12);
 assign p_18_13 = p_18_15 & p_14_13;
 assign g_18_13 = g_18_15 | (p_18_15 & g_14_13);
 assign p_18_14 = p_18_15 & p_14_14;
 assign g_18_14 = g_18_15 | (p_18_15 & g_14_14);
 assign p_18_15 = p_18_17 & p_16_15;
 assign g_18_15 = g_18_17 | (p_18_17 & g_16_15);
 assign p_18_16 = p_18_17 & p_16_16;
 assign g_18_16 = g_18_17 | (p_18_17 & g_16_16);
 assign p_18_17 = p_18_18 & p_17_17;
 assign g_18_17 = g_18_18 | (p_18_18 & g_17_17);
 assign sum[18] = p_18_18^ g_17_0;
 assign p_19_0 = p_19_4 & p_3_0;
 assign g_19_0 = g_19_4 | (p_19_4 & g_3_0);
 assign p_19_1 = p_19_4 & p_3_1;
 assign g_19_1 = g_19_4 | (p_19_4 & g_3_1);
 assign p_19_2 = p_19_4 & p_3_2;
 assign g_19_2 = g_19_4 | (p_19_4 & g_3_2);
 assign p_19_3 = p_19_4 & p_3_3;
 assign g_19_3 = g_19_4 | (p_19_4 & g_3_3);
 assign p_19_4 = p_19_12 & p_11_4;
 assign g_19_4 = g_19_12 | (p_19_12 & g_11_4);
 assign p_19_5 = p_19_12 & p_11_5;
 assign g_19_5 = g_19_12 | (p_19_12 & g_11_5);
 assign p_19_6 = p_19_12 & p_11_6;
 assign g_19_6 = g_19_12 | (p_19_12 & g_11_6);
 assign p_19_7 = p_19_12 & p_11_7;
 assign g_19_7 = g_19_12 | (p_19_12 & g_11_7);
 assign p_19_8 = p_19_12 & p_11_8;
 assign g_19_8 = g_19_12 | (p_19_12 & g_11_8);
 assign p_19_9 = p_19_12 & p_11_9;
 assign g_19_9 = g_19_12 | (p_19_12 & g_11_9);
 assign p_19_10 = p_19_12 & p_11_10;
 assign g_19_10 = g_19_12 | (p_19_12 & g_11_10);
 assign p_19_11 = p_19_12 & p_11_11;
 assign g_19_11 = g_19_12 | (p_19_12 & g_11_11);
 assign p_19_12 = p_19_16 & p_15_12;
 assign g_19_12 = g_19_16 | (p_19_16 & g_15_12);
 assign p_19_13 = p_19_16 & p_15_13;
 assign g_19_13 = g_19_16 | (p_19_16 & g_15_13);
 assign p_19_14 = p_19_16 & p_15_14;
 assign g_19_14 = g_19_16 | (p_19_16 & g_15_14);
 assign p_19_15 = p_19_16 & p_15_15;
 assign g_19_15 = g_19_16 | (p_19_16 & g_15_15);
 assign p_19_16 = p_19_18 & p_17_16;
 assign g_19_16 = g_19_18 | (p_19_18 & g_17_16);
 assign p_19_17 = p_19_18 & p_17_17;
 assign g_19_17 = g_19_18 | (p_19_18 & g_17_17);
 assign p_19_18 = p_19_19 & p_18_18;
 assign g_19_18 = g_19_19 | (p_19_19 & g_18_18);
 assign sum[19] = p_19_19^ g_18_0;
 assign p_20_0 = p_20_5 & p_4_0;
 assign g_20_0 = g_20_5 | (p_20_5 & g_4_0);
 assign p_20_1 = p_20_5 & p_4_1;
 assign g_20_1 = g_20_5 | (p_20_5 & g_4_1);
 assign p_20_2 = p_20_5 & p_4_2;
 assign g_20_2 = g_20_5 | (p_20_5 & g_4_2);
 assign p_20_3 = p_20_5 & p_4_3;
 assign g_20_3 = g_20_5 | (p_20_5 & g_4_3);
 assign p_20_4 = p_20_5 & p_4_4;
 assign g_20_4 = g_20_5 | (p_20_5 & g_4_4);
 assign p_20_5 = p_20_13 & p_12_5;
 assign g_20_5 = g_20_13 | (p_20_13 & g_12_5);
 assign p_20_6 = p_20_13 & p_12_6;
 assign g_20_6 = g_20_13 | (p_20_13 & g_12_6);
 assign p_20_7 = p_20_13 & p_12_7;
 assign g_20_7 = g_20_13 | (p_20_13 & g_12_7);
 assign p_20_8 = p_20_13 & p_12_8;
 assign g_20_8 = g_20_13 | (p_20_13 & g_12_8);
 assign p_20_9 = p_20_13 & p_12_9;
 assign g_20_9 = g_20_13 | (p_20_13 & g_12_9);
 assign p_20_10 = p_20_13 & p_12_10;
 assign g_20_10 = g_20_13 | (p_20_13 & g_12_10);
 assign p_20_11 = p_20_13 & p_12_11;
 assign g_20_11 = g_20_13 | (p_20_13 & g_12_11);
 assign p_20_12 = p_20_13 & p_12_12;
 assign g_20_12 = g_20_13 | (p_20_13 & g_12_12);
 assign p_20_13 = p_20_17 & p_16_13;
 assign g_20_13 = g_20_17 | (p_20_17 & g_16_13);
 assign p_20_14 = p_20_17 & p_16_14;
 assign g_20_14 = g_20_17 | (p_20_17 & g_16_14);
 assign p_20_15 = p_20_17 & p_16_15;
 assign g_20_15 = g_20_17 | (p_20_17 & g_16_15);
 assign p_20_16 = p_20_17 & p_16_16;
 assign g_20_16 = g_20_17 | (p_20_17 & g_16_16);
 assign p_20_17 = p_20_19 & p_18_17;
 assign g_20_17 = g_20_19 | (p_20_19 & g_18_17);
 assign p_20_18 = p_20_19 & p_18_18;
 assign g_20_18 = g_20_19 | (p_20_19 & g_18_18);
 assign p_20_19 = p_20_20 & p_19_19;
 assign g_20_19 = g_20_20 | (p_20_20 & g_19_19);
 assign sum[20] = p_20_20^ g_19_0;
 assign p_21_0 = p_21_6 & p_5_0;
 assign g_21_0 = g_21_6 | (p_21_6 & g_5_0);
 assign p_21_1 = p_21_6 & p_5_1;
 assign g_21_1 = g_21_6 | (p_21_6 & g_5_1);
 assign p_21_2 = p_21_6 & p_5_2;
 assign g_21_2 = g_21_6 | (p_21_6 & g_5_2);
 assign p_21_3 = p_21_6 & p_5_3;
 assign g_21_3 = g_21_6 | (p_21_6 & g_5_3);
 assign p_21_4 = p_21_6 & p_5_4;
 assign g_21_4 = g_21_6 | (p_21_6 & g_5_4);
 assign p_21_5 = p_21_6 & p_5_5;
 assign g_21_5 = g_21_6 | (p_21_6 & g_5_5);
 assign p_21_6 = p_21_14 & p_13_6;
 assign g_21_6 = g_21_14 | (p_21_14 & g_13_6);
 assign p_21_7 = p_21_14 & p_13_7;
 assign g_21_7 = g_21_14 | (p_21_14 & g_13_7);
 assign p_21_8 = p_21_14 & p_13_8;
 assign g_21_8 = g_21_14 | (p_21_14 & g_13_8);
 assign p_21_9 = p_21_14 & p_13_9;
 assign g_21_9 = g_21_14 | (p_21_14 & g_13_9);
 assign p_21_10 = p_21_14 & p_13_10;
 assign g_21_10 = g_21_14 | (p_21_14 & g_13_10);
 assign p_21_11 = p_21_14 & p_13_11;
 assign g_21_11 = g_21_14 | (p_21_14 & g_13_11);
 assign p_21_12 = p_21_14 & p_13_12;
 assign g_21_12 = g_21_14 | (p_21_14 & g_13_12);
 assign p_21_13 = p_21_14 & p_13_13;
 assign g_21_13 = g_21_14 | (p_21_14 & g_13_13);
 assign p_21_14 = p_21_18 & p_17_14;
 assign g_21_14 = g_21_18 | (p_21_18 & g_17_14);
 assign p_21_15 = p_21_18 & p_17_15;
 assign g_21_15 = g_21_18 | (p_21_18 & g_17_15);
 assign p_21_16 = p_21_18 & p_17_16;
 assign g_21_16 = g_21_18 | (p_21_18 & g_17_16);
 assign p_21_17 = p_21_18 & p_17_17;
 assign g_21_17 = g_21_18 | (p_21_18 & g_17_17);
 assign p_21_18 = p_21_20 & p_19_18;
 assign g_21_18 = g_21_20 | (p_21_20 & g_19_18);
 assign p_21_19 = p_21_20 & p_19_19;
 assign g_21_19 = g_21_20 | (p_21_20 & g_19_19);
 assign p_21_20 = p_21_21 & p_20_20;
 assign g_21_20 = g_21_21 | (p_21_21 & g_20_20);
 assign sum[21] = p_21_21^ g_20_0;
 assign p_22_0 = p_22_7 & p_6_0;
 assign g_22_0 = g_22_7 | (p_22_7 & g_6_0);
 assign p_22_1 = p_22_7 & p_6_1;
 assign g_22_1 = g_22_7 | (p_22_7 & g_6_1);
 assign p_22_2 = p_22_7 & p_6_2;
 assign g_22_2 = g_22_7 | (p_22_7 & g_6_2);
 assign p_22_3 = p_22_7 & p_6_3;
 assign g_22_3 = g_22_7 | (p_22_7 & g_6_3);
 assign p_22_4 = p_22_7 & p_6_4;
 assign g_22_4 = g_22_7 | (p_22_7 & g_6_4);
 assign p_22_5 = p_22_7 & p_6_5;
 assign g_22_5 = g_22_7 | (p_22_7 & g_6_5);
 assign p_22_6 = p_22_7 & p_6_6;
 assign g_22_6 = g_22_7 | (p_22_7 & g_6_6);
 assign p_22_7 = p_22_15 & p_14_7;
 assign g_22_7 = g_22_15 | (p_22_15 & g_14_7);
 assign p_22_8 = p_22_15 & p_14_8;
 assign g_22_8 = g_22_15 | (p_22_15 & g_14_8);
 assign p_22_9 = p_22_15 & p_14_9;
 assign g_22_9 = g_22_15 | (p_22_15 & g_14_9);
 assign p_22_10 = p_22_15 & p_14_10;
 assign g_22_10 = g_22_15 | (p_22_15 & g_14_10);
 assign p_22_11 = p_22_15 & p_14_11;
 assign g_22_11 = g_22_15 | (p_22_15 & g_14_11);
 assign p_22_12 = p_22_15 & p_14_12;
 assign g_22_12 = g_22_15 | (p_22_15 & g_14_12);
 assign p_22_13 = p_22_15 & p_14_13;
 assign g_22_13 = g_22_15 | (p_22_15 & g_14_13);
 assign p_22_14 = p_22_15 & p_14_14;
 assign g_22_14 = g_22_15 | (p_22_15 & g_14_14);
 assign p_22_15 = p_22_19 & p_18_15;
 assign g_22_15 = g_22_19 | (p_22_19 & g_18_15);
 assign p_22_16 = p_22_19 & p_18_16;
 assign g_22_16 = g_22_19 | (p_22_19 & g_18_16);
 assign p_22_17 = p_22_19 & p_18_17;
 assign g_22_17 = g_22_19 | (p_22_19 & g_18_17);
 assign p_22_18 = p_22_19 & p_18_18;
 assign g_22_18 = g_22_19 | (p_22_19 & g_18_18);
 assign p_22_19 = p_22_21 & p_20_19;
 assign g_22_19 = g_22_21 | (p_22_21 & g_20_19);
 assign p_22_20 = p_22_21 & p_20_20;
 assign g_22_20 = g_22_21 | (p_22_21 & g_20_20);
 assign p_22_21 = p_22_22 & p_21_21;
 assign g_22_21 = g_22_22 | (p_22_22 & g_21_21);
 assign sum[22] = p_22_22^ g_21_0;
 assign p_23_0 = p_23_8 & p_7_0;
 assign g_23_0 = g_23_8 | (p_23_8 & g_7_0);
 assign p_23_1 = p_23_8 & p_7_1;
 assign g_23_1 = g_23_8 | (p_23_8 & g_7_1);
 assign p_23_2 = p_23_8 & p_7_2;
 assign g_23_2 = g_23_8 | (p_23_8 & g_7_2);
 assign p_23_3 = p_23_8 & p_7_3;
 assign g_23_3 = g_23_8 | (p_23_8 & g_7_3);
 assign p_23_4 = p_23_8 & p_7_4;
 assign g_23_4 = g_23_8 | (p_23_8 & g_7_4);
 assign p_23_5 = p_23_8 & p_7_5;
 assign g_23_5 = g_23_8 | (p_23_8 & g_7_5);
 assign p_23_6 = p_23_8 & p_7_6;
 assign g_23_6 = g_23_8 | (p_23_8 & g_7_6);
 assign p_23_7 = p_23_8 & p_7_7;
 assign g_23_7 = g_23_8 | (p_23_8 & g_7_7);
 assign p_23_8 = p_23_16 & p_15_8;
 assign g_23_8 = g_23_16 | (p_23_16 & g_15_8);
 assign p_23_9 = p_23_16 & p_15_9;
 assign g_23_9 = g_23_16 | (p_23_16 & g_15_9);
 assign p_23_10 = p_23_16 & p_15_10;
 assign g_23_10 = g_23_16 | (p_23_16 & g_15_10);
 assign p_23_11 = p_23_16 & p_15_11;
 assign g_23_11 = g_23_16 | (p_23_16 & g_15_11);
 assign p_23_12 = p_23_16 & p_15_12;
 assign g_23_12 = g_23_16 | (p_23_16 & g_15_12);
 assign p_23_13 = p_23_16 & p_15_13;
 assign g_23_13 = g_23_16 | (p_23_16 & g_15_13);
 assign p_23_14 = p_23_16 & p_15_14;
 assign g_23_14 = g_23_16 | (p_23_16 & g_15_14);
 assign p_23_15 = p_23_16 & p_15_15;
 assign g_23_15 = g_23_16 | (p_23_16 & g_15_15);
 assign p_23_16 = p_23_20 & p_19_16;
 assign g_23_16 = g_23_20 | (p_23_20 & g_19_16);
 assign p_23_17 = p_23_20 & p_19_17;
 assign g_23_17 = g_23_20 | (p_23_20 & g_19_17);
 assign p_23_18 = p_23_20 & p_19_18;
 assign g_23_18 = g_23_20 | (p_23_20 & g_19_18);
 assign p_23_19 = p_23_20 & p_19_19;
 assign g_23_19 = g_23_20 | (p_23_20 & g_19_19);
 assign p_23_20 = p_23_22 & p_21_20;
 assign g_23_20 = g_23_22 | (p_23_22 & g_21_20);
 assign p_23_21 = p_23_22 & p_21_21;
 assign g_23_21 = g_23_22 | (p_23_22 & g_21_21);
 assign p_23_22 = p_23_23 & p_22_22;
 assign g_23_22 = g_23_23 | (p_23_23 & g_22_22);
 assign sum[23] = p_23_23^ g_22_0;
 assign p_24_0 = p_24_9 & p_8_0;
 assign g_24_0 = g_24_9 | (p_24_9 & g_8_0);
 assign p_24_1 = p_24_9 & p_8_1;
 assign g_24_1 = g_24_9 | (p_24_9 & g_8_1);
 assign p_24_2 = p_24_9 & p_8_2;
 assign g_24_2 = g_24_9 | (p_24_9 & g_8_2);
 assign p_24_3 = p_24_9 & p_8_3;
 assign g_24_3 = g_24_9 | (p_24_9 & g_8_3);
 assign p_24_4 = p_24_9 & p_8_4;
 assign g_24_4 = g_24_9 | (p_24_9 & g_8_4);
 assign p_24_5 = p_24_9 & p_8_5;
 assign g_24_5 = g_24_9 | (p_24_9 & g_8_5);
 assign p_24_6 = p_24_9 & p_8_6;
 assign g_24_6 = g_24_9 | (p_24_9 & g_8_6);
 assign p_24_7 = p_24_9 & p_8_7;
 assign g_24_7 = g_24_9 | (p_24_9 & g_8_7);
 assign p_24_8 = p_24_9 & p_8_8;
 assign g_24_8 = g_24_9 | (p_24_9 & g_8_8);
 assign p_24_9 = p_24_17 & p_16_9;
 assign g_24_9 = g_24_17 | (p_24_17 & g_16_9);
 assign p_24_10 = p_24_17 & p_16_10;
 assign g_24_10 = g_24_17 | (p_24_17 & g_16_10);
 assign p_24_11 = p_24_17 & p_16_11;
 assign g_24_11 = g_24_17 | (p_24_17 & g_16_11);
 assign p_24_12 = p_24_17 & p_16_12;
 assign g_24_12 = g_24_17 | (p_24_17 & g_16_12);
 assign p_24_13 = p_24_17 & p_16_13;
 assign g_24_13 = g_24_17 | (p_24_17 & g_16_13);
 assign p_24_14 = p_24_17 & p_16_14;
 assign g_24_14 = g_24_17 | (p_24_17 & g_16_14);
 assign p_24_15 = p_24_17 & p_16_15;
 assign g_24_15 = g_24_17 | (p_24_17 & g_16_15);
 assign p_24_16 = p_24_17 & p_16_16;
 assign g_24_16 = g_24_17 | (p_24_17 & g_16_16);
 assign p_24_17 = p_24_21 & p_20_17;
 assign g_24_17 = g_24_21 | (p_24_21 & g_20_17);
 assign p_24_18 = p_24_21 & p_20_18;
 assign g_24_18 = g_24_21 | (p_24_21 & g_20_18);
 assign p_24_19 = p_24_21 & p_20_19;
 assign g_24_19 = g_24_21 | (p_24_21 & g_20_19);
 assign p_24_20 = p_24_21 & p_20_20;
 assign g_24_20 = g_24_21 | (p_24_21 & g_20_20);
 assign p_24_21 = p_24_23 & p_22_21;
 assign g_24_21 = g_24_23 | (p_24_23 & g_22_21);
 assign p_24_22 = p_24_23 & p_22_22;
 assign g_24_22 = g_24_23 | (p_24_23 & g_22_22);
 assign p_24_23 = p_24_24 & p_23_23;
 assign g_24_23 = g_24_24 | (p_24_24 & g_23_23);
 assign sum[24] = p_24_24^ g_23_0;
 assign p_25_0 = p_25_10 & p_9_0;
 assign g_25_0 = g_25_10 | (p_25_10 & g_9_0);
 assign p_25_1 = p_25_10 & p_9_1;
 assign g_25_1 = g_25_10 | (p_25_10 & g_9_1);
 assign p_25_2 = p_25_10 & p_9_2;
 assign g_25_2 = g_25_10 | (p_25_10 & g_9_2);
 assign p_25_3 = p_25_10 & p_9_3;
 assign g_25_3 = g_25_10 | (p_25_10 & g_9_3);
 assign p_25_4 = p_25_10 & p_9_4;
 assign g_25_4 = g_25_10 | (p_25_10 & g_9_4);
 assign p_25_5 = p_25_10 & p_9_5;
 assign g_25_5 = g_25_10 | (p_25_10 & g_9_5);
 assign p_25_6 = p_25_10 & p_9_6;
 assign g_25_6 = g_25_10 | (p_25_10 & g_9_6);
 assign p_25_7 = p_25_10 & p_9_7;
 assign g_25_7 = g_25_10 | (p_25_10 & g_9_7);
 assign p_25_8 = p_25_10 & p_9_8;
 assign g_25_8 = g_25_10 | (p_25_10 & g_9_8);
 assign p_25_9 = p_25_10 & p_9_9;
 assign g_25_9 = g_25_10 | (p_25_10 & g_9_9);
 assign p_25_10 = p_25_18 & p_17_10;
 assign g_25_10 = g_25_18 | (p_25_18 & g_17_10);
 assign p_25_11 = p_25_18 & p_17_11;
 assign g_25_11 = g_25_18 | (p_25_18 & g_17_11);
 assign p_25_12 = p_25_18 & p_17_12;
 assign g_25_12 = g_25_18 | (p_25_18 & g_17_12);
 assign p_25_13 = p_25_18 & p_17_13;
 assign g_25_13 = g_25_18 | (p_25_18 & g_17_13);
 assign p_25_14 = p_25_18 & p_17_14;
 assign g_25_14 = g_25_18 | (p_25_18 & g_17_14);
 assign p_25_15 = p_25_18 & p_17_15;
 assign g_25_15 = g_25_18 | (p_25_18 & g_17_15);
 assign p_25_16 = p_25_18 & p_17_16;
 assign g_25_16 = g_25_18 | (p_25_18 & g_17_16);
 assign p_25_17 = p_25_18 & p_17_17;
 assign g_25_17 = g_25_18 | (p_25_18 & g_17_17);
 assign p_25_18 = p_25_22 & p_21_18;
 assign g_25_18 = g_25_22 | (p_25_22 & g_21_18);
 assign p_25_19 = p_25_22 & p_21_19;
 assign g_25_19 = g_25_22 | (p_25_22 & g_21_19);
 assign p_25_20 = p_25_22 & p_21_20;
 assign g_25_20 = g_25_22 | (p_25_22 & g_21_20);
 assign p_25_21 = p_25_22 & p_21_21;
 assign g_25_21 = g_25_22 | (p_25_22 & g_21_21);
 assign p_25_22 = p_25_24 & p_23_22;
 assign g_25_22 = g_25_24 | (p_25_24 & g_23_22);
 assign p_25_23 = p_25_24 & p_23_23;
 assign g_25_23 = g_25_24 | (p_25_24 & g_23_23);
 assign p_25_24 = p_25_25 & p_24_24;
 assign g_25_24 = g_25_25 | (p_25_25 & g_24_24);
 assign sum[25] = p_25_25^ g_24_0;
 assign p_26_0 = p_26_11 & p_10_0;
 assign g_26_0 = g_26_11 | (p_26_11 & g_10_0);
 assign p_26_1 = p_26_11 & p_10_1;
 assign g_26_1 = g_26_11 | (p_26_11 & g_10_1);
 assign p_26_2 = p_26_11 & p_10_2;
 assign g_26_2 = g_26_11 | (p_26_11 & g_10_2);
 assign p_26_3 = p_26_11 & p_10_3;
 assign g_26_3 = g_26_11 | (p_26_11 & g_10_3);
 assign p_26_4 = p_26_11 & p_10_4;
 assign g_26_4 = g_26_11 | (p_26_11 & g_10_4);
 assign p_26_5 = p_26_11 & p_10_5;
 assign g_26_5 = g_26_11 | (p_26_11 & g_10_5);
 assign p_26_6 = p_26_11 & p_10_6;
 assign g_26_6 = g_26_11 | (p_26_11 & g_10_6);
 assign p_26_7 = p_26_11 & p_10_7;
 assign g_26_7 = g_26_11 | (p_26_11 & g_10_7);
 assign p_26_8 = p_26_11 & p_10_8;
 assign g_26_8 = g_26_11 | (p_26_11 & g_10_8);
 assign p_26_9 = p_26_11 & p_10_9;
 assign g_26_9 = g_26_11 | (p_26_11 & g_10_9);
 assign p_26_10 = p_26_11 & p_10_10;
 assign g_26_10 = g_26_11 | (p_26_11 & g_10_10);
 assign p_26_11 = p_26_19 & p_18_11;
 assign g_26_11 = g_26_19 | (p_26_19 & g_18_11);
 assign p_26_12 = p_26_19 & p_18_12;
 assign g_26_12 = g_26_19 | (p_26_19 & g_18_12);
 assign p_26_13 = p_26_19 & p_18_13;
 assign g_26_13 = g_26_19 | (p_26_19 & g_18_13);
 assign p_26_14 = p_26_19 & p_18_14;
 assign g_26_14 = g_26_19 | (p_26_19 & g_18_14);
 assign p_26_15 = p_26_19 & p_18_15;
 assign g_26_15 = g_26_19 | (p_26_19 & g_18_15);
 assign p_26_16 = p_26_19 & p_18_16;
 assign g_26_16 = g_26_19 | (p_26_19 & g_18_16);
 assign p_26_17 = p_26_19 & p_18_17;
 assign g_26_17 = g_26_19 | (p_26_19 & g_18_17);
 assign p_26_18 = p_26_19 & p_18_18;
 assign g_26_18 = g_26_19 | (p_26_19 & g_18_18);
 assign p_26_19 = p_26_23 & p_22_19;
 assign g_26_19 = g_26_23 | (p_26_23 & g_22_19);
 assign p_26_20 = p_26_23 & p_22_20;
 assign g_26_20 = g_26_23 | (p_26_23 & g_22_20);
 assign p_26_21 = p_26_23 & p_22_21;
 assign g_26_21 = g_26_23 | (p_26_23 & g_22_21);
 assign p_26_22 = p_26_23 & p_22_22;
 assign g_26_22 = g_26_23 | (p_26_23 & g_22_22);
 assign p_26_23 = p_26_25 & p_24_23;
 assign g_26_23 = g_26_25 | (p_26_25 & g_24_23);
 assign p_26_24 = p_26_25 & p_24_24;
 assign g_26_24 = g_26_25 | (p_26_25 & g_24_24);
 assign p_26_25 = p_26_26 & p_25_25;
 assign g_26_25 = g_26_26 | (p_26_26 & g_25_25);
 assign sum[26] = p_26_26^ g_25_0;
 assign p_27_0 = p_27_12 & p_11_0;
 assign g_27_0 = g_27_12 | (p_27_12 & g_11_0);
 assign p_27_1 = p_27_12 & p_11_1;
 assign g_27_1 = g_27_12 | (p_27_12 & g_11_1);
 assign p_27_2 = p_27_12 & p_11_2;
 assign g_27_2 = g_27_12 | (p_27_12 & g_11_2);
 assign p_27_3 = p_27_12 & p_11_3;
 assign g_27_3 = g_27_12 | (p_27_12 & g_11_3);
 assign p_27_4 = p_27_12 & p_11_4;
 assign g_27_4 = g_27_12 | (p_27_12 & g_11_4);
 assign p_27_5 = p_27_12 & p_11_5;
 assign g_27_5 = g_27_12 | (p_27_12 & g_11_5);
 assign p_27_6 = p_27_12 & p_11_6;
 assign g_27_6 = g_27_12 | (p_27_12 & g_11_6);
 assign p_27_7 = p_27_12 & p_11_7;
 assign g_27_7 = g_27_12 | (p_27_12 & g_11_7);
 assign p_27_8 = p_27_12 & p_11_8;
 assign g_27_8 = g_27_12 | (p_27_12 & g_11_8);
 assign p_27_9 = p_27_12 & p_11_9;
 assign g_27_9 = g_27_12 | (p_27_12 & g_11_9);
 assign p_27_10 = p_27_12 & p_11_10;
 assign g_27_10 = g_27_12 | (p_27_12 & g_11_10);
 assign p_27_11 = p_27_12 & p_11_11;
 assign g_27_11 = g_27_12 | (p_27_12 & g_11_11);
 assign p_27_12 = p_27_20 & p_19_12;
 assign g_27_12 = g_27_20 | (p_27_20 & g_19_12);
 assign p_27_13 = p_27_20 & p_19_13;
 assign g_27_13 = g_27_20 | (p_27_20 & g_19_13);
 assign p_27_14 = p_27_20 & p_19_14;
 assign g_27_14 = g_27_20 | (p_27_20 & g_19_14);
 assign p_27_15 = p_27_20 & p_19_15;
 assign g_27_15 = g_27_20 | (p_27_20 & g_19_15);
 assign p_27_16 = p_27_20 & p_19_16;
 assign g_27_16 = g_27_20 | (p_27_20 & g_19_16);
 assign p_27_17 = p_27_20 & p_19_17;
 assign g_27_17 = g_27_20 | (p_27_20 & g_19_17);
 assign p_27_18 = p_27_20 & p_19_18;
 assign g_27_18 = g_27_20 | (p_27_20 & g_19_18);
 assign p_27_19 = p_27_20 & p_19_19;
 assign g_27_19 = g_27_20 | (p_27_20 & g_19_19);
 assign p_27_20 = p_27_24 & p_23_20;
 assign g_27_20 = g_27_24 | (p_27_24 & g_23_20);
 assign p_27_21 = p_27_24 & p_23_21;
 assign g_27_21 = g_27_24 | (p_27_24 & g_23_21);
 assign p_27_22 = p_27_24 & p_23_22;
 assign g_27_22 = g_27_24 | (p_27_24 & g_23_22);
 assign p_27_23 = p_27_24 & p_23_23;
 assign g_27_23 = g_27_24 | (p_27_24 & g_23_23);
 assign p_27_24 = p_27_26 & p_25_24;
 assign g_27_24 = g_27_26 | (p_27_26 & g_25_24);
 assign p_27_25 = p_27_26 & p_25_25;
 assign g_27_25 = g_27_26 | (p_27_26 & g_25_25);
 assign p_27_26 = p_27_27 & p_26_26;
 assign g_27_26 = g_27_27 | (p_27_27 & g_26_26);
 assign sum[27] = p_27_27^ g_26_0;
 assign p_28_0 = p_28_13 & p_12_0;
 assign g_28_0 = g_28_13 | (p_28_13 & g_12_0);
 assign p_28_1 = p_28_13 & p_12_1;
 assign g_28_1 = g_28_13 | (p_28_13 & g_12_1);
 assign p_28_2 = p_28_13 & p_12_2;
 assign g_28_2 = g_28_13 | (p_28_13 & g_12_2);
 assign p_28_3 = p_28_13 & p_12_3;
 assign g_28_3 = g_28_13 | (p_28_13 & g_12_3);
 assign p_28_4 = p_28_13 & p_12_4;
 assign g_28_4 = g_28_13 | (p_28_13 & g_12_4);
 assign p_28_5 = p_28_13 & p_12_5;
 assign g_28_5 = g_28_13 | (p_28_13 & g_12_5);
 assign p_28_6 = p_28_13 & p_12_6;
 assign g_28_6 = g_28_13 | (p_28_13 & g_12_6);
 assign p_28_7 = p_28_13 & p_12_7;
 assign g_28_7 = g_28_13 | (p_28_13 & g_12_7);
 assign p_28_8 = p_28_13 & p_12_8;
 assign g_28_8 = g_28_13 | (p_28_13 & g_12_8);
 assign p_28_9 = p_28_13 & p_12_9;
 assign g_28_9 = g_28_13 | (p_28_13 & g_12_9);
 assign p_28_10 = p_28_13 & p_12_10;
 assign g_28_10 = g_28_13 | (p_28_13 & g_12_10);
 assign p_28_11 = p_28_13 & p_12_11;
 assign g_28_11 = g_28_13 | (p_28_13 & g_12_11);
 assign p_28_12 = p_28_13 & p_12_12;
 assign g_28_12 = g_28_13 | (p_28_13 & g_12_12);
 assign p_28_13 = p_28_21 & p_20_13;
 assign g_28_13 = g_28_21 | (p_28_21 & g_20_13);
 assign p_28_14 = p_28_21 & p_20_14;
 assign g_28_14 = g_28_21 | (p_28_21 & g_20_14);
 assign p_28_15 = p_28_21 & p_20_15;
 assign g_28_15 = g_28_21 | (p_28_21 & g_20_15);
 assign p_28_16 = p_28_21 & p_20_16;
 assign g_28_16 = g_28_21 | (p_28_21 & g_20_16);
 assign p_28_17 = p_28_21 & p_20_17;
 assign g_28_17 = g_28_21 | (p_28_21 & g_20_17);
 assign p_28_18 = p_28_21 & p_20_18;
 assign g_28_18 = g_28_21 | (p_28_21 & g_20_18);
 assign p_28_19 = p_28_21 & p_20_19;
 assign g_28_19 = g_28_21 | (p_28_21 & g_20_19);
 assign p_28_20 = p_28_21 & p_20_20;
 assign g_28_20 = g_28_21 | (p_28_21 & g_20_20);
 assign p_28_21 = p_28_25 & p_24_21;
 assign g_28_21 = g_28_25 | (p_28_25 & g_24_21);
 assign p_28_22 = p_28_25 & p_24_22;
 assign g_28_22 = g_28_25 | (p_28_25 & g_24_22);
 assign p_28_23 = p_28_25 & p_24_23;
 assign g_28_23 = g_28_25 | (p_28_25 & g_24_23);
 assign p_28_24 = p_28_25 & p_24_24;
 assign g_28_24 = g_28_25 | (p_28_25 & g_24_24);
 assign p_28_25 = p_28_27 & p_26_25;
 assign g_28_25 = g_28_27 | (p_28_27 & g_26_25);
 assign p_28_26 = p_28_27 & p_26_26;
 assign g_28_26 = g_28_27 | (p_28_27 & g_26_26);
 assign p_28_27 = p_28_28 & p_27_27;
 assign g_28_27 = g_28_28 | (p_28_28 & g_27_27);
 assign sum[28] = p_28_28^ g_27_0;
 assign p_29_0 = p_29_14 & p_13_0;
 assign g_29_0 = g_29_14 | (p_29_14 & g_13_0);
 assign p_29_1 = p_29_14 & p_13_1;
 assign g_29_1 = g_29_14 | (p_29_14 & g_13_1);
 assign p_29_2 = p_29_14 & p_13_2;
 assign g_29_2 = g_29_14 | (p_29_14 & g_13_2);
 assign p_29_3 = p_29_14 & p_13_3;
 assign g_29_3 = g_29_14 | (p_29_14 & g_13_3);
 assign p_29_4 = p_29_14 & p_13_4;
 assign g_29_4 = g_29_14 | (p_29_14 & g_13_4);
 assign p_29_5 = p_29_14 & p_13_5;
 assign g_29_5 = g_29_14 | (p_29_14 & g_13_5);
 assign p_29_6 = p_29_14 & p_13_6;
 assign g_29_6 = g_29_14 | (p_29_14 & g_13_6);
 assign p_29_7 = p_29_14 & p_13_7;
 assign g_29_7 = g_29_14 | (p_29_14 & g_13_7);
 assign p_29_8 = p_29_14 & p_13_8;
 assign g_29_8 = g_29_14 | (p_29_14 & g_13_8);
 assign p_29_9 = p_29_14 & p_13_9;
 assign g_29_9 = g_29_14 | (p_29_14 & g_13_9);
 assign p_29_10 = p_29_14 & p_13_10;
 assign g_29_10 = g_29_14 | (p_29_14 & g_13_10);
 assign p_29_11 = p_29_14 & p_13_11;
 assign g_29_11 = g_29_14 | (p_29_14 & g_13_11);
 assign p_29_12 = p_29_14 & p_13_12;
 assign g_29_12 = g_29_14 | (p_29_14 & g_13_12);
 assign p_29_13 = p_29_14 & p_13_13;
 assign g_29_13 = g_29_14 | (p_29_14 & g_13_13);
 assign p_29_14 = p_29_22 & p_21_14;
 assign g_29_14 = g_29_22 | (p_29_22 & g_21_14);
 assign p_29_15 = p_29_22 & p_21_15;
 assign g_29_15 = g_29_22 | (p_29_22 & g_21_15);
 assign p_29_16 = p_29_22 & p_21_16;
 assign g_29_16 = g_29_22 | (p_29_22 & g_21_16);
 assign p_29_17 = p_29_22 & p_21_17;
 assign g_29_17 = g_29_22 | (p_29_22 & g_21_17);
 assign p_29_18 = p_29_22 & p_21_18;
 assign g_29_18 = g_29_22 | (p_29_22 & g_21_18);
 assign p_29_19 = p_29_22 & p_21_19;
 assign g_29_19 = g_29_22 | (p_29_22 & g_21_19);
 assign p_29_20 = p_29_22 & p_21_20;
 assign g_29_20 = g_29_22 | (p_29_22 & g_21_20);
 assign p_29_21 = p_29_22 & p_21_21;
 assign g_29_21 = g_29_22 | (p_29_22 & g_21_21);
 assign p_29_22 = p_29_26 & p_25_22;
 assign g_29_22 = g_29_26 | (p_29_26 & g_25_22);
 assign p_29_23 = p_29_26 & p_25_23;
 assign g_29_23 = g_29_26 | (p_29_26 & g_25_23);
 assign p_29_24 = p_29_26 & p_25_24;
 assign g_29_24 = g_29_26 | (p_29_26 & g_25_24);
 assign p_29_25 = p_29_26 & p_25_25;
 assign g_29_25 = g_29_26 | (p_29_26 & g_25_25);
 assign p_29_26 = p_29_28 & p_27_26;
 assign g_29_26 = g_29_28 | (p_29_28 & g_27_26);
 assign p_29_27 = p_29_28 & p_27_27;
 assign g_29_27 = g_29_28 | (p_29_28 & g_27_27);
 assign p_29_28 = p_29_29 & p_28_28;
 assign g_29_28 = g_29_29 | (p_29_29 & g_28_28);
 assign sum[29] = p_29_29^ g_28_0;
 assign p_30_0 = p_30_15 & p_14_0;
 assign g_30_0 = g_30_15 | (p_30_15 & g_14_0);
 assign p_30_1 = p_30_15 & p_14_1;
 assign g_30_1 = g_30_15 | (p_30_15 & g_14_1);
 assign p_30_2 = p_30_15 & p_14_2;
 assign g_30_2 = g_30_15 | (p_30_15 & g_14_2);
 assign p_30_3 = p_30_15 & p_14_3;
 assign g_30_3 = g_30_15 | (p_30_15 & g_14_3);
 assign p_30_4 = p_30_15 & p_14_4;
 assign g_30_4 = g_30_15 | (p_30_15 & g_14_4);
 assign p_30_5 = p_30_15 & p_14_5;
 assign g_30_5 = g_30_15 | (p_30_15 & g_14_5);
 assign p_30_6 = p_30_15 & p_14_6;
 assign g_30_6 = g_30_15 | (p_30_15 & g_14_6);
 assign p_30_7 = p_30_15 & p_14_7;
 assign g_30_7 = g_30_15 | (p_30_15 & g_14_7);
 assign p_30_8 = p_30_15 & p_14_8;
 assign g_30_8 = g_30_15 | (p_30_15 & g_14_8);
 assign p_30_9 = p_30_15 & p_14_9;
 assign g_30_9 = g_30_15 | (p_30_15 & g_14_9);
 assign p_30_10 = p_30_15 & p_14_10;
 assign g_30_10 = g_30_15 | (p_30_15 & g_14_10);
 assign p_30_11 = p_30_15 & p_14_11;
 assign g_30_11 = g_30_15 | (p_30_15 & g_14_11);
 assign p_30_12 = p_30_15 & p_14_12;
 assign g_30_12 = g_30_15 | (p_30_15 & g_14_12);
 assign p_30_13 = p_30_15 & p_14_13;
 assign g_30_13 = g_30_15 | (p_30_15 & g_14_13);
 assign p_30_14 = p_30_15 & p_14_14;
 assign g_30_14 = g_30_15 | (p_30_15 & g_14_14);
 assign p_30_15 = p_30_23 & p_22_15;
 assign g_30_15 = g_30_23 | (p_30_23 & g_22_15);
 assign p_30_16 = p_30_23 & p_22_16;
 assign g_30_16 = g_30_23 | (p_30_23 & g_22_16);
 assign p_30_17 = p_30_23 & p_22_17;
 assign g_30_17 = g_30_23 | (p_30_23 & g_22_17);
 assign p_30_18 = p_30_23 & p_22_18;
 assign g_30_18 = g_30_23 | (p_30_23 & g_22_18);
 assign p_30_19 = p_30_23 & p_22_19;
 assign g_30_19 = g_30_23 | (p_30_23 & g_22_19);
 assign p_30_20 = p_30_23 & p_22_20;
 assign g_30_20 = g_30_23 | (p_30_23 & g_22_20);
 assign p_30_21 = p_30_23 & p_22_21;
 assign g_30_21 = g_30_23 | (p_30_23 & g_22_21);
 assign p_30_22 = p_30_23 & p_22_22;
 assign g_30_22 = g_30_23 | (p_30_23 & g_22_22);
 assign p_30_23 = p_30_27 & p_26_23;
 assign g_30_23 = g_30_27 | (p_30_27 & g_26_23);
 assign p_30_24 = p_30_27 & p_26_24;
 assign g_30_24 = g_30_27 | (p_30_27 & g_26_24);
 assign p_30_25 = p_30_27 & p_26_25;
 assign g_30_25 = g_30_27 | (p_30_27 & g_26_25);
 assign p_30_26 = p_30_27 & p_26_26;
 assign g_30_26 = g_30_27 | (p_30_27 & g_26_26);
 assign p_30_27 = p_30_29 & p_28_27;
 assign g_30_27 = g_30_29 | (p_30_29 & g_28_27);
 assign p_30_28 = p_30_29 & p_28_28;
 assign g_30_28 = g_30_29 | (p_30_29 & g_28_28);
 assign p_30_29 = p_30_30 & p_29_29;
 assign g_30_29 = g_30_30 | (p_30_30 & g_29_29);
 assign sum[30] = p_30_30^ g_29_0;
 assign cout = g_30_0;
endmodule
