module MG_FA(
  input a,
  input b,
  input cin,
  output sum,
  output cout
);

  assign sum = (a ^ b) ^ cin;
  assign cout = (a & b) | (b & cin) | (a & cin);
endmodule
module MG_HA(
  input a,
  input b,
  output sum,
  output cout
);

  assign sum = a ^ b;
  assign cout = a & b;
endmodule
module mult32u_booth4_sklansky(
  input [31:0] multiplicand,
  input [31:0] multiplier,
  output [63:0] product
);

  wire be_2x_0_0;
  wire be_2x_0_1;
  wire be_2x_0_10;
  wire be_2x_0_11;
  wire be_2x_0_12;
  wire be_2x_0_13;
  wire be_2x_0_14;
  wire be_2x_0_15;
  wire be_2x_0_16;
  wire be_2x_0_17;
  wire be_2x_0_18;
  wire be_2x_0_19;
  wire be_2x_0_2;
  wire be_2x_0_20;
  wire be_2x_0_21;
  wire be_2x_0_22;
  wire be_2x_0_23;
  wire be_2x_0_24;
  wire be_2x_0_25;
  wire be_2x_0_26;
  wire be_2x_0_27;
  wire be_2x_0_28;
  wire be_2x_0_29;
  wire be_2x_0_3;
  wire be_2x_0_30;
  wire be_2x_0_31;
  wire be_2x_0_32;
  wire be_2x_0_33;
  wire be_2x_0_4;
  wire be_2x_0_5;
  wire be_2x_0_6;
  wire be_2x_0_7;
  wire be_2x_0_8;
  wire be_2x_0_9;
  wire be_2x_10_0;
  wire be_2x_10_1;
  wire be_2x_10_10;
  wire be_2x_10_11;
  wire be_2x_10_12;
  wire be_2x_10_13;
  wire be_2x_10_14;
  wire be_2x_10_15;
  wire be_2x_10_16;
  wire be_2x_10_17;
  wire be_2x_10_18;
  wire be_2x_10_19;
  wire be_2x_10_2;
  wire be_2x_10_20;
  wire be_2x_10_21;
  wire be_2x_10_22;
  wire be_2x_10_23;
  wire be_2x_10_24;
  wire be_2x_10_25;
  wire be_2x_10_26;
  wire be_2x_10_27;
  wire be_2x_10_28;
  wire be_2x_10_29;
  wire be_2x_10_3;
  wire be_2x_10_30;
  wire be_2x_10_31;
  wire be_2x_10_32;
  wire be_2x_10_33;
  wire be_2x_10_4;
  wire be_2x_10_5;
  wire be_2x_10_6;
  wire be_2x_10_7;
  wire be_2x_10_8;
  wire be_2x_10_9;
  wire be_2x_11_0;
  wire be_2x_11_1;
  wire be_2x_11_10;
  wire be_2x_11_11;
  wire be_2x_11_12;
  wire be_2x_11_13;
  wire be_2x_11_14;
  wire be_2x_11_15;
  wire be_2x_11_16;
  wire be_2x_11_17;
  wire be_2x_11_18;
  wire be_2x_11_19;
  wire be_2x_11_2;
  wire be_2x_11_20;
  wire be_2x_11_21;
  wire be_2x_11_22;
  wire be_2x_11_23;
  wire be_2x_11_24;
  wire be_2x_11_25;
  wire be_2x_11_26;
  wire be_2x_11_27;
  wire be_2x_11_28;
  wire be_2x_11_29;
  wire be_2x_11_3;
  wire be_2x_11_30;
  wire be_2x_11_31;
  wire be_2x_11_32;
  wire be_2x_11_33;
  wire be_2x_11_4;
  wire be_2x_11_5;
  wire be_2x_11_6;
  wire be_2x_11_7;
  wire be_2x_11_8;
  wire be_2x_11_9;
  wire be_2x_12_0;
  wire be_2x_12_1;
  wire be_2x_12_10;
  wire be_2x_12_11;
  wire be_2x_12_12;
  wire be_2x_12_13;
  wire be_2x_12_14;
  wire be_2x_12_15;
  wire be_2x_12_16;
  wire be_2x_12_17;
  wire be_2x_12_18;
  wire be_2x_12_19;
  wire be_2x_12_2;
  wire be_2x_12_20;
  wire be_2x_12_21;
  wire be_2x_12_22;
  wire be_2x_12_23;
  wire be_2x_12_24;
  wire be_2x_12_25;
  wire be_2x_12_26;
  wire be_2x_12_27;
  wire be_2x_12_28;
  wire be_2x_12_29;
  wire be_2x_12_3;
  wire be_2x_12_30;
  wire be_2x_12_31;
  wire be_2x_12_32;
  wire be_2x_12_33;
  wire be_2x_12_4;
  wire be_2x_12_5;
  wire be_2x_12_6;
  wire be_2x_12_7;
  wire be_2x_12_8;
  wire be_2x_12_9;
  wire be_2x_13_0;
  wire be_2x_13_1;
  wire be_2x_13_10;
  wire be_2x_13_11;
  wire be_2x_13_12;
  wire be_2x_13_13;
  wire be_2x_13_14;
  wire be_2x_13_15;
  wire be_2x_13_16;
  wire be_2x_13_17;
  wire be_2x_13_18;
  wire be_2x_13_19;
  wire be_2x_13_2;
  wire be_2x_13_20;
  wire be_2x_13_21;
  wire be_2x_13_22;
  wire be_2x_13_23;
  wire be_2x_13_24;
  wire be_2x_13_25;
  wire be_2x_13_26;
  wire be_2x_13_27;
  wire be_2x_13_28;
  wire be_2x_13_29;
  wire be_2x_13_3;
  wire be_2x_13_30;
  wire be_2x_13_31;
  wire be_2x_13_32;
  wire be_2x_13_33;
  wire be_2x_13_4;
  wire be_2x_13_5;
  wire be_2x_13_6;
  wire be_2x_13_7;
  wire be_2x_13_8;
  wire be_2x_13_9;
  wire be_2x_14_0;
  wire be_2x_14_1;
  wire be_2x_14_10;
  wire be_2x_14_11;
  wire be_2x_14_12;
  wire be_2x_14_13;
  wire be_2x_14_14;
  wire be_2x_14_15;
  wire be_2x_14_16;
  wire be_2x_14_17;
  wire be_2x_14_18;
  wire be_2x_14_19;
  wire be_2x_14_2;
  wire be_2x_14_20;
  wire be_2x_14_21;
  wire be_2x_14_22;
  wire be_2x_14_23;
  wire be_2x_14_24;
  wire be_2x_14_25;
  wire be_2x_14_26;
  wire be_2x_14_27;
  wire be_2x_14_28;
  wire be_2x_14_29;
  wire be_2x_14_3;
  wire be_2x_14_30;
  wire be_2x_14_31;
  wire be_2x_14_32;
  wire be_2x_14_33;
  wire be_2x_14_4;
  wire be_2x_14_5;
  wire be_2x_14_6;
  wire be_2x_14_7;
  wire be_2x_14_8;
  wire be_2x_14_9;
  wire be_2x_15_0;
  wire be_2x_15_1;
  wire be_2x_15_10;
  wire be_2x_15_11;
  wire be_2x_15_12;
  wire be_2x_15_13;
  wire be_2x_15_14;
  wire be_2x_15_15;
  wire be_2x_15_16;
  wire be_2x_15_17;
  wire be_2x_15_18;
  wire be_2x_15_19;
  wire be_2x_15_2;
  wire be_2x_15_20;
  wire be_2x_15_21;
  wire be_2x_15_22;
  wire be_2x_15_23;
  wire be_2x_15_24;
  wire be_2x_15_25;
  wire be_2x_15_26;
  wire be_2x_15_27;
  wire be_2x_15_28;
  wire be_2x_15_29;
  wire be_2x_15_3;
  wire be_2x_15_30;
  wire be_2x_15_31;
  wire be_2x_15_32;
  wire be_2x_15_33;
  wire be_2x_15_4;
  wire be_2x_15_5;
  wire be_2x_15_6;
  wire be_2x_15_7;
  wire be_2x_15_8;
  wire be_2x_15_9;
  wire be_2x_16_0;
  wire be_2x_16_1;
  wire be_2x_16_10;
  wire be_2x_16_11;
  wire be_2x_16_12;
  wire be_2x_16_13;
  wire be_2x_16_14;
  wire be_2x_16_15;
  wire be_2x_16_16;
  wire be_2x_16_17;
  wire be_2x_16_18;
  wire be_2x_16_19;
  wire be_2x_16_2;
  wire be_2x_16_20;
  wire be_2x_16_21;
  wire be_2x_16_22;
  wire be_2x_16_23;
  wire be_2x_16_24;
  wire be_2x_16_25;
  wire be_2x_16_26;
  wire be_2x_16_27;
  wire be_2x_16_28;
  wire be_2x_16_29;
  wire be_2x_16_3;
  wire be_2x_16_30;
  wire be_2x_16_31;
  wire be_2x_16_4;
  wire be_2x_16_5;
  wire be_2x_16_6;
  wire be_2x_16_7;
  wire be_2x_16_8;
  wire be_2x_16_9;
  wire be_2x_1_0;
  wire be_2x_1_1;
  wire be_2x_1_10;
  wire be_2x_1_11;
  wire be_2x_1_12;
  wire be_2x_1_13;
  wire be_2x_1_14;
  wire be_2x_1_15;
  wire be_2x_1_16;
  wire be_2x_1_17;
  wire be_2x_1_18;
  wire be_2x_1_19;
  wire be_2x_1_2;
  wire be_2x_1_20;
  wire be_2x_1_21;
  wire be_2x_1_22;
  wire be_2x_1_23;
  wire be_2x_1_24;
  wire be_2x_1_25;
  wire be_2x_1_26;
  wire be_2x_1_27;
  wire be_2x_1_28;
  wire be_2x_1_29;
  wire be_2x_1_3;
  wire be_2x_1_30;
  wire be_2x_1_31;
  wire be_2x_1_32;
  wire be_2x_1_33;
  wire be_2x_1_4;
  wire be_2x_1_5;
  wire be_2x_1_6;
  wire be_2x_1_7;
  wire be_2x_1_8;
  wire be_2x_1_9;
  wire be_2x_2_0;
  wire be_2x_2_1;
  wire be_2x_2_10;
  wire be_2x_2_11;
  wire be_2x_2_12;
  wire be_2x_2_13;
  wire be_2x_2_14;
  wire be_2x_2_15;
  wire be_2x_2_16;
  wire be_2x_2_17;
  wire be_2x_2_18;
  wire be_2x_2_19;
  wire be_2x_2_2;
  wire be_2x_2_20;
  wire be_2x_2_21;
  wire be_2x_2_22;
  wire be_2x_2_23;
  wire be_2x_2_24;
  wire be_2x_2_25;
  wire be_2x_2_26;
  wire be_2x_2_27;
  wire be_2x_2_28;
  wire be_2x_2_29;
  wire be_2x_2_3;
  wire be_2x_2_30;
  wire be_2x_2_31;
  wire be_2x_2_32;
  wire be_2x_2_33;
  wire be_2x_2_4;
  wire be_2x_2_5;
  wire be_2x_2_6;
  wire be_2x_2_7;
  wire be_2x_2_8;
  wire be_2x_2_9;
  wire be_2x_3_0;
  wire be_2x_3_1;
  wire be_2x_3_10;
  wire be_2x_3_11;
  wire be_2x_3_12;
  wire be_2x_3_13;
  wire be_2x_3_14;
  wire be_2x_3_15;
  wire be_2x_3_16;
  wire be_2x_3_17;
  wire be_2x_3_18;
  wire be_2x_3_19;
  wire be_2x_3_2;
  wire be_2x_3_20;
  wire be_2x_3_21;
  wire be_2x_3_22;
  wire be_2x_3_23;
  wire be_2x_3_24;
  wire be_2x_3_25;
  wire be_2x_3_26;
  wire be_2x_3_27;
  wire be_2x_3_28;
  wire be_2x_3_29;
  wire be_2x_3_3;
  wire be_2x_3_30;
  wire be_2x_3_31;
  wire be_2x_3_32;
  wire be_2x_3_33;
  wire be_2x_3_4;
  wire be_2x_3_5;
  wire be_2x_3_6;
  wire be_2x_3_7;
  wire be_2x_3_8;
  wire be_2x_3_9;
  wire be_2x_4_0;
  wire be_2x_4_1;
  wire be_2x_4_10;
  wire be_2x_4_11;
  wire be_2x_4_12;
  wire be_2x_4_13;
  wire be_2x_4_14;
  wire be_2x_4_15;
  wire be_2x_4_16;
  wire be_2x_4_17;
  wire be_2x_4_18;
  wire be_2x_4_19;
  wire be_2x_4_2;
  wire be_2x_4_20;
  wire be_2x_4_21;
  wire be_2x_4_22;
  wire be_2x_4_23;
  wire be_2x_4_24;
  wire be_2x_4_25;
  wire be_2x_4_26;
  wire be_2x_4_27;
  wire be_2x_4_28;
  wire be_2x_4_29;
  wire be_2x_4_3;
  wire be_2x_4_30;
  wire be_2x_4_31;
  wire be_2x_4_32;
  wire be_2x_4_33;
  wire be_2x_4_4;
  wire be_2x_4_5;
  wire be_2x_4_6;
  wire be_2x_4_7;
  wire be_2x_4_8;
  wire be_2x_4_9;
  wire be_2x_5_0;
  wire be_2x_5_1;
  wire be_2x_5_10;
  wire be_2x_5_11;
  wire be_2x_5_12;
  wire be_2x_5_13;
  wire be_2x_5_14;
  wire be_2x_5_15;
  wire be_2x_5_16;
  wire be_2x_5_17;
  wire be_2x_5_18;
  wire be_2x_5_19;
  wire be_2x_5_2;
  wire be_2x_5_20;
  wire be_2x_5_21;
  wire be_2x_5_22;
  wire be_2x_5_23;
  wire be_2x_5_24;
  wire be_2x_5_25;
  wire be_2x_5_26;
  wire be_2x_5_27;
  wire be_2x_5_28;
  wire be_2x_5_29;
  wire be_2x_5_3;
  wire be_2x_5_30;
  wire be_2x_5_31;
  wire be_2x_5_32;
  wire be_2x_5_33;
  wire be_2x_5_4;
  wire be_2x_5_5;
  wire be_2x_5_6;
  wire be_2x_5_7;
  wire be_2x_5_8;
  wire be_2x_5_9;
  wire be_2x_6_0;
  wire be_2x_6_1;
  wire be_2x_6_10;
  wire be_2x_6_11;
  wire be_2x_6_12;
  wire be_2x_6_13;
  wire be_2x_6_14;
  wire be_2x_6_15;
  wire be_2x_6_16;
  wire be_2x_6_17;
  wire be_2x_6_18;
  wire be_2x_6_19;
  wire be_2x_6_2;
  wire be_2x_6_20;
  wire be_2x_6_21;
  wire be_2x_6_22;
  wire be_2x_6_23;
  wire be_2x_6_24;
  wire be_2x_6_25;
  wire be_2x_6_26;
  wire be_2x_6_27;
  wire be_2x_6_28;
  wire be_2x_6_29;
  wire be_2x_6_3;
  wire be_2x_6_30;
  wire be_2x_6_31;
  wire be_2x_6_32;
  wire be_2x_6_33;
  wire be_2x_6_4;
  wire be_2x_6_5;
  wire be_2x_6_6;
  wire be_2x_6_7;
  wire be_2x_6_8;
  wire be_2x_6_9;
  wire be_2x_7_0;
  wire be_2x_7_1;
  wire be_2x_7_10;
  wire be_2x_7_11;
  wire be_2x_7_12;
  wire be_2x_7_13;
  wire be_2x_7_14;
  wire be_2x_7_15;
  wire be_2x_7_16;
  wire be_2x_7_17;
  wire be_2x_7_18;
  wire be_2x_7_19;
  wire be_2x_7_2;
  wire be_2x_7_20;
  wire be_2x_7_21;
  wire be_2x_7_22;
  wire be_2x_7_23;
  wire be_2x_7_24;
  wire be_2x_7_25;
  wire be_2x_7_26;
  wire be_2x_7_27;
  wire be_2x_7_28;
  wire be_2x_7_29;
  wire be_2x_7_3;
  wire be_2x_7_30;
  wire be_2x_7_31;
  wire be_2x_7_32;
  wire be_2x_7_33;
  wire be_2x_7_4;
  wire be_2x_7_5;
  wire be_2x_7_6;
  wire be_2x_7_7;
  wire be_2x_7_8;
  wire be_2x_7_9;
  wire be_2x_8_0;
  wire be_2x_8_1;
  wire be_2x_8_10;
  wire be_2x_8_11;
  wire be_2x_8_12;
  wire be_2x_8_13;
  wire be_2x_8_14;
  wire be_2x_8_15;
  wire be_2x_8_16;
  wire be_2x_8_17;
  wire be_2x_8_18;
  wire be_2x_8_19;
  wire be_2x_8_2;
  wire be_2x_8_20;
  wire be_2x_8_21;
  wire be_2x_8_22;
  wire be_2x_8_23;
  wire be_2x_8_24;
  wire be_2x_8_25;
  wire be_2x_8_26;
  wire be_2x_8_27;
  wire be_2x_8_28;
  wire be_2x_8_29;
  wire be_2x_8_3;
  wire be_2x_8_30;
  wire be_2x_8_31;
  wire be_2x_8_32;
  wire be_2x_8_33;
  wire be_2x_8_4;
  wire be_2x_8_5;
  wire be_2x_8_6;
  wire be_2x_8_7;
  wire be_2x_8_8;
  wire be_2x_8_9;
  wire be_2x_9_0;
  wire be_2x_9_1;
  wire be_2x_9_10;
  wire be_2x_9_11;
  wire be_2x_9_12;
  wire be_2x_9_13;
  wire be_2x_9_14;
  wire be_2x_9_15;
  wire be_2x_9_16;
  wire be_2x_9_17;
  wire be_2x_9_18;
  wire be_2x_9_19;
  wire be_2x_9_2;
  wire be_2x_9_20;
  wire be_2x_9_21;
  wire be_2x_9_22;
  wire be_2x_9_23;
  wire be_2x_9_24;
  wire be_2x_9_25;
  wire be_2x_9_26;
  wire be_2x_9_27;
  wire be_2x_9_28;
  wire be_2x_9_29;
  wire be_2x_9_3;
  wire be_2x_9_30;
  wire be_2x_9_31;
  wire be_2x_9_32;
  wire be_2x_9_33;
  wire be_2x_9_4;
  wire be_2x_9_5;
  wire be_2x_9_6;
  wire be_2x_9_7;
  wire be_2x_9_8;
  wire be_2x_9_9;
  wire be_c_0;
  wire be_c_1;
  wire be_c_10;
  wire be_c_11;
  wire be_c_12;
  wire be_c_13;
  wire be_c_14;
  wire be_c_15;
  wire be_c_16;
  wire be_c_2;
  wire be_c_3;
  wire be_c_4;
  wire be_c_5;
  wire be_c_6;
  wire be_c_7;
  wire be_c_8;
  wire be_c_9;
  wire be_d_0;
  wire be_d_1;
  wire be_d_10;
  wire be_d_11;
  wire be_d_12;
  wire be_d_13;
  wire be_d_14;
  wire be_d_15;
  wire be_d_16;
  wire be_d_2;
  wire be_d_3;
  wire be_d_4;
  wire be_d_5;
  wire be_d_6;
  wire be_d_7;
  wire be_d_8;
  wire be_d_9;
  wire be_neg_0;
  wire be_neg_1;
  wire be_neg_10;
  wire be_neg_11;
  wire be_neg_12;
  wire be_neg_13;
  wire be_neg_14;
  wire be_neg_15;
  wire be_neg_16;
  wire be_neg_2;
  wire be_neg_3;
  wire be_neg_4;
  wire be_neg_5;
  wire be_neg_6;
  wire be_neg_7;
  wire be_neg_8;
  wire be_neg_9;
  wire be_s1_0;
  wire be_s1_1;
  wire be_s1_10;
  wire be_s1_11;
  wire be_s1_12;
  wire be_s1_13;
  wire be_s1_14;
  wire be_s1_15;
  wire be_s1_16;
  wire be_s1_2;
  wire be_s1_3;
  wire be_s1_4;
  wire be_s1_5;
  wire be_s1_6;
  wire be_s1_7;
  wire be_s1_8;
  wire be_s1_9;
  wire be_s2_0;
  wire be_s2_1;
  wire be_s2_10;
  wire be_s2_11;
  wire be_s2_12;
  wire be_s2_13;
  wire be_s2_14;
  wire be_s2_15;
  wire be_s2_16;
  wire be_s2_2;
  wire be_s2_3;
  wire be_s2_4;
  wire be_s2_5;
  wire be_s2_6;
  wire be_s2_7;
  wire be_s2_8;
  wire be_s2_9;
  wire be_s2_a_0;
  wire be_s2_a_1;
  wire be_s2_a_10;
  wire be_s2_a_11;
  wire be_s2_a_12;
  wire be_s2_a_13;
  wire be_s2_a_14;
  wire be_s2_a_15;
  wire be_s2_a_16;
  wire be_s2_a_2;
  wire be_s2_a_3;
  wire be_s2_a_4;
  wire be_s2_a_5;
  wire be_s2_a_6;
  wire be_s2_a_7;
  wire be_s2_a_8;
  wire be_s2_a_9;
  wire be_s2_b_0;
  wire be_s2_b_1;
  wire be_s2_b_10;
  wire be_s2_b_11;
  wire be_s2_b_12;
  wire be_s2_b_13;
  wire be_s2_b_14;
  wire be_s2_b_15;
  wire be_s2_b_16;
  wire be_s2_b_2;
  wire be_s2_b_3;
  wire be_s2_b_4;
  wire be_s2_b_5;
  wire be_s2_b_6;
  wire be_s2_b_7;
  wire be_s2_b_8;
  wire be_s2_b_9;
  wire be_x_0_0;
  wire be_x_0_1;
  wire be_x_0_10;
  wire be_x_0_11;
  wire be_x_0_12;
  wire be_x_0_13;
  wire be_x_0_14;
  wire be_x_0_15;
  wire be_x_0_16;
  wire be_x_0_17;
  wire be_x_0_18;
  wire be_x_0_19;
  wire be_x_0_2;
  wire be_x_0_20;
  wire be_x_0_21;
  wire be_x_0_22;
  wire be_x_0_23;
  wire be_x_0_24;
  wire be_x_0_25;
  wire be_x_0_26;
  wire be_x_0_27;
  wire be_x_0_28;
  wire be_x_0_29;
  wire be_x_0_3;
  wire be_x_0_30;
  wire be_x_0_31;
  wire be_x_0_32;
  wire be_x_0_33;
  wire be_x_0_4;
  wire be_x_0_5;
  wire be_x_0_6;
  wire be_x_0_7;
  wire be_x_0_8;
  wire be_x_0_9;
  wire be_x_10_0;
  wire be_x_10_1;
  wire be_x_10_10;
  wire be_x_10_11;
  wire be_x_10_12;
  wire be_x_10_13;
  wire be_x_10_14;
  wire be_x_10_15;
  wire be_x_10_16;
  wire be_x_10_17;
  wire be_x_10_18;
  wire be_x_10_19;
  wire be_x_10_2;
  wire be_x_10_20;
  wire be_x_10_21;
  wire be_x_10_22;
  wire be_x_10_23;
  wire be_x_10_24;
  wire be_x_10_25;
  wire be_x_10_26;
  wire be_x_10_27;
  wire be_x_10_28;
  wire be_x_10_29;
  wire be_x_10_3;
  wire be_x_10_30;
  wire be_x_10_31;
  wire be_x_10_32;
  wire be_x_10_33;
  wire be_x_10_4;
  wire be_x_10_5;
  wire be_x_10_6;
  wire be_x_10_7;
  wire be_x_10_8;
  wire be_x_10_9;
  wire be_x_11_0;
  wire be_x_11_1;
  wire be_x_11_10;
  wire be_x_11_11;
  wire be_x_11_12;
  wire be_x_11_13;
  wire be_x_11_14;
  wire be_x_11_15;
  wire be_x_11_16;
  wire be_x_11_17;
  wire be_x_11_18;
  wire be_x_11_19;
  wire be_x_11_2;
  wire be_x_11_20;
  wire be_x_11_21;
  wire be_x_11_22;
  wire be_x_11_23;
  wire be_x_11_24;
  wire be_x_11_25;
  wire be_x_11_26;
  wire be_x_11_27;
  wire be_x_11_28;
  wire be_x_11_29;
  wire be_x_11_3;
  wire be_x_11_30;
  wire be_x_11_31;
  wire be_x_11_32;
  wire be_x_11_33;
  wire be_x_11_4;
  wire be_x_11_5;
  wire be_x_11_6;
  wire be_x_11_7;
  wire be_x_11_8;
  wire be_x_11_9;
  wire be_x_12_0;
  wire be_x_12_1;
  wire be_x_12_10;
  wire be_x_12_11;
  wire be_x_12_12;
  wire be_x_12_13;
  wire be_x_12_14;
  wire be_x_12_15;
  wire be_x_12_16;
  wire be_x_12_17;
  wire be_x_12_18;
  wire be_x_12_19;
  wire be_x_12_2;
  wire be_x_12_20;
  wire be_x_12_21;
  wire be_x_12_22;
  wire be_x_12_23;
  wire be_x_12_24;
  wire be_x_12_25;
  wire be_x_12_26;
  wire be_x_12_27;
  wire be_x_12_28;
  wire be_x_12_29;
  wire be_x_12_3;
  wire be_x_12_30;
  wire be_x_12_31;
  wire be_x_12_32;
  wire be_x_12_33;
  wire be_x_12_4;
  wire be_x_12_5;
  wire be_x_12_6;
  wire be_x_12_7;
  wire be_x_12_8;
  wire be_x_12_9;
  wire be_x_13_0;
  wire be_x_13_1;
  wire be_x_13_10;
  wire be_x_13_11;
  wire be_x_13_12;
  wire be_x_13_13;
  wire be_x_13_14;
  wire be_x_13_15;
  wire be_x_13_16;
  wire be_x_13_17;
  wire be_x_13_18;
  wire be_x_13_19;
  wire be_x_13_2;
  wire be_x_13_20;
  wire be_x_13_21;
  wire be_x_13_22;
  wire be_x_13_23;
  wire be_x_13_24;
  wire be_x_13_25;
  wire be_x_13_26;
  wire be_x_13_27;
  wire be_x_13_28;
  wire be_x_13_29;
  wire be_x_13_3;
  wire be_x_13_30;
  wire be_x_13_31;
  wire be_x_13_32;
  wire be_x_13_33;
  wire be_x_13_4;
  wire be_x_13_5;
  wire be_x_13_6;
  wire be_x_13_7;
  wire be_x_13_8;
  wire be_x_13_9;
  wire be_x_14_0;
  wire be_x_14_1;
  wire be_x_14_10;
  wire be_x_14_11;
  wire be_x_14_12;
  wire be_x_14_13;
  wire be_x_14_14;
  wire be_x_14_15;
  wire be_x_14_16;
  wire be_x_14_17;
  wire be_x_14_18;
  wire be_x_14_19;
  wire be_x_14_2;
  wire be_x_14_20;
  wire be_x_14_21;
  wire be_x_14_22;
  wire be_x_14_23;
  wire be_x_14_24;
  wire be_x_14_25;
  wire be_x_14_26;
  wire be_x_14_27;
  wire be_x_14_28;
  wire be_x_14_29;
  wire be_x_14_3;
  wire be_x_14_30;
  wire be_x_14_31;
  wire be_x_14_32;
  wire be_x_14_33;
  wire be_x_14_4;
  wire be_x_14_5;
  wire be_x_14_6;
  wire be_x_14_7;
  wire be_x_14_8;
  wire be_x_14_9;
  wire be_x_15_0;
  wire be_x_15_1;
  wire be_x_15_10;
  wire be_x_15_11;
  wire be_x_15_12;
  wire be_x_15_13;
  wire be_x_15_14;
  wire be_x_15_15;
  wire be_x_15_16;
  wire be_x_15_17;
  wire be_x_15_18;
  wire be_x_15_19;
  wire be_x_15_2;
  wire be_x_15_20;
  wire be_x_15_21;
  wire be_x_15_22;
  wire be_x_15_23;
  wire be_x_15_24;
  wire be_x_15_25;
  wire be_x_15_26;
  wire be_x_15_27;
  wire be_x_15_28;
  wire be_x_15_29;
  wire be_x_15_3;
  wire be_x_15_30;
  wire be_x_15_31;
  wire be_x_15_32;
  wire be_x_15_33;
  wire be_x_15_4;
  wire be_x_15_5;
  wire be_x_15_6;
  wire be_x_15_7;
  wire be_x_15_8;
  wire be_x_15_9;
  wire be_x_16_0;
  wire be_x_16_1;
  wire be_x_16_10;
  wire be_x_16_11;
  wire be_x_16_12;
  wire be_x_16_13;
  wire be_x_16_14;
  wire be_x_16_15;
  wire be_x_16_16;
  wire be_x_16_17;
  wire be_x_16_18;
  wire be_x_16_19;
  wire be_x_16_2;
  wire be_x_16_20;
  wire be_x_16_21;
  wire be_x_16_22;
  wire be_x_16_23;
  wire be_x_16_24;
  wire be_x_16_25;
  wire be_x_16_26;
  wire be_x_16_27;
  wire be_x_16_28;
  wire be_x_16_29;
  wire be_x_16_3;
  wire be_x_16_30;
  wire be_x_16_31;
  wire be_x_16_4;
  wire be_x_16_5;
  wire be_x_16_6;
  wire be_x_16_7;
  wire be_x_16_8;
  wire be_x_16_9;
  wire be_x_1_0;
  wire be_x_1_1;
  wire be_x_1_10;
  wire be_x_1_11;
  wire be_x_1_12;
  wire be_x_1_13;
  wire be_x_1_14;
  wire be_x_1_15;
  wire be_x_1_16;
  wire be_x_1_17;
  wire be_x_1_18;
  wire be_x_1_19;
  wire be_x_1_2;
  wire be_x_1_20;
  wire be_x_1_21;
  wire be_x_1_22;
  wire be_x_1_23;
  wire be_x_1_24;
  wire be_x_1_25;
  wire be_x_1_26;
  wire be_x_1_27;
  wire be_x_1_28;
  wire be_x_1_29;
  wire be_x_1_3;
  wire be_x_1_30;
  wire be_x_1_31;
  wire be_x_1_32;
  wire be_x_1_33;
  wire be_x_1_4;
  wire be_x_1_5;
  wire be_x_1_6;
  wire be_x_1_7;
  wire be_x_1_8;
  wire be_x_1_9;
  wire be_x_2_0;
  wire be_x_2_1;
  wire be_x_2_10;
  wire be_x_2_11;
  wire be_x_2_12;
  wire be_x_2_13;
  wire be_x_2_14;
  wire be_x_2_15;
  wire be_x_2_16;
  wire be_x_2_17;
  wire be_x_2_18;
  wire be_x_2_19;
  wire be_x_2_2;
  wire be_x_2_20;
  wire be_x_2_21;
  wire be_x_2_22;
  wire be_x_2_23;
  wire be_x_2_24;
  wire be_x_2_25;
  wire be_x_2_26;
  wire be_x_2_27;
  wire be_x_2_28;
  wire be_x_2_29;
  wire be_x_2_3;
  wire be_x_2_30;
  wire be_x_2_31;
  wire be_x_2_32;
  wire be_x_2_33;
  wire be_x_2_4;
  wire be_x_2_5;
  wire be_x_2_6;
  wire be_x_2_7;
  wire be_x_2_8;
  wire be_x_2_9;
  wire be_x_3_0;
  wire be_x_3_1;
  wire be_x_3_10;
  wire be_x_3_11;
  wire be_x_3_12;
  wire be_x_3_13;
  wire be_x_3_14;
  wire be_x_3_15;
  wire be_x_3_16;
  wire be_x_3_17;
  wire be_x_3_18;
  wire be_x_3_19;
  wire be_x_3_2;
  wire be_x_3_20;
  wire be_x_3_21;
  wire be_x_3_22;
  wire be_x_3_23;
  wire be_x_3_24;
  wire be_x_3_25;
  wire be_x_3_26;
  wire be_x_3_27;
  wire be_x_3_28;
  wire be_x_3_29;
  wire be_x_3_3;
  wire be_x_3_30;
  wire be_x_3_31;
  wire be_x_3_32;
  wire be_x_3_33;
  wire be_x_3_4;
  wire be_x_3_5;
  wire be_x_3_6;
  wire be_x_3_7;
  wire be_x_3_8;
  wire be_x_3_9;
  wire be_x_4_0;
  wire be_x_4_1;
  wire be_x_4_10;
  wire be_x_4_11;
  wire be_x_4_12;
  wire be_x_4_13;
  wire be_x_4_14;
  wire be_x_4_15;
  wire be_x_4_16;
  wire be_x_4_17;
  wire be_x_4_18;
  wire be_x_4_19;
  wire be_x_4_2;
  wire be_x_4_20;
  wire be_x_4_21;
  wire be_x_4_22;
  wire be_x_4_23;
  wire be_x_4_24;
  wire be_x_4_25;
  wire be_x_4_26;
  wire be_x_4_27;
  wire be_x_4_28;
  wire be_x_4_29;
  wire be_x_4_3;
  wire be_x_4_30;
  wire be_x_4_31;
  wire be_x_4_32;
  wire be_x_4_33;
  wire be_x_4_4;
  wire be_x_4_5;
  wire be_x_4_6;
  wire be_x_4_7;
  wire be_x_4_8;
  wire be_x_4_9;
  wire be_x_5_0;
  wire be_x_5_1;
  wire be_x_5_10;
  wire be_x_5_11;
  wire be_x_5_12;
  wire be_x_5_13;
  wire be_x_5_14;
  wire be_x_5_15;
  wire be_x_5_16;
  wire be_x_5_17;
  wire be_x_5_18;
  wire be_x_5_19;
  wire be_x_5_2;
  wire be_x_5_20;
  wire be_x_5_21;
  wire be_x_5_22;
  wire be_x_5_23;
  wire be_x_5_24;
  wire be_x_5_25;
  wire be_x_5_26;
  wire be_x_5_27;
  wire be_x_5_28;
  wire be_x_5_29;
  wire be_x_5_3;
  wire be_x_5_30;
  wire be_x_5_31;
  wire be_x_5_32;
  wire be_x_5_33;
  wire be_x_5_4;
  wire be_x_5_5;
  wire be_x_5_6;
  wire be_x_5_7;
  wire be_x_5_8;
  wire be_x_5_9;
  wire be_x_6_0;
  wire be_x_6_1;
  wire be_x_6_10;
  wire be_x_6_11;
  wire be_x_6_12;
  wire be_x_6_13;
  wire be_x_6_14;
  wire be_x_6_15;
  wire be_x_6_16;
  wire be_x_6_17;
  wire be_x_6_18;
  wire be_x_6_19;
  wire be_x_6_2;
  wire be_x_6_20;
  wire be_x_6_21;
  wire be_x_6_22;
  wire be_x_6_23;
  wire be_x_6_24;
  wire be_x_6_25;
  wire be_x_6_26;
  wire be_x_6_27;
  wire be_x_6_28;
  wire be_x_6_29;
  wire be_x_6_3;
  wire be_x_6_30;
  wire be_x_6_31;
  wire be_x_6_32;
  wire be_x_6_33;
  wire be_x_6_4;
  wire be_x_6_5;
  wire be_x_6_6;
  wire be_x_6_7;
  wire be_x_6_8;
  wire be_x_6_9;
  wire be_x_7_0;
  wire be_x_7_1;
  wire be_x_7_10;
  wire be_x_7_11;
  wire be_x_7_12;
  wire be_x_7_13;
  wire be_x_7_14;
  wire be_x_7_15;
  wire be_x_7_16;
  wire be_x_7_17;
  wire be_x_7_18;
  wire be_x_7_19;
  wire be_x_7_2;
  wire be_x_7_20;
  wire be_x_7_21;
  wire be_x_7_22;
  wire be_x_7_23;
  wire be_x_7_24;
  wire be_x_7_25;
  wire be_x_7_26;
  wire be_x_7_27;
  wire be_x_7_28;
  wire be_x_7_29;
  wire be_x_7_3;
  wire be_x_7_30;
  wire be_x_7_31;
  wire be_x_7_32;
  wire be_x_7_33;
  wire be_x_7_4;
  wire be_x_7_5;
  wire be_x_7_6;
  wire be_x_7_7;
  wire be_x_7_8;
  wire be_x_7_9;
  wire be_x_8_0;
  wire be_x_8_1;
  wire be_x_8_10;
  wire be_x_8_11;
  wire be_x_8_12;
  wire be_x_8_13;
  wire be_x_8_14;
  wire be_x_8_15;
  wire be_x_8_16;
  wire be_x_8_17;
  wire be_x_8_18;
  wire be_x_8_19;
  wire be_x_8_2;
  wire be_x_8_20;
  wire be_x_8_21;
  wire be_x_8_22;
  wire be_x_8_23;
  wire be_x_8_24;
  wire be_x_8_25;
  wire be_x_8_26;
  wire be_x_8_27;
  wire be_x_8_28;
  wire be_x_8_29;
  wire be_x_8_3;
  wire be_x_8_30;
  wire be_x_8_31;
  wire be_x_8_32;
  wire be_x_8_33;
  wire be_x_8_4;
  wire be_x_8_5;
  wire be_x_8_6;
  wire be_x_8_7;
  wire be_x_8_8;
  wire be_x_8_9;
  wire be_x_9_0;
  wire be_x_9_1;
  wire be_x_9_10;
  wire be_x_9_11;
  wire be_x_9_12;
  wire be_x_9_13;
  wire be_x_9_14;
  wire be_x_9_15;
  wire be_x_9_16;
  wire be_x_9_17;
  wire be_x_9_18;
  wire be_x_9_19;
  wire be_x_9_2;
  wire be_x_9_20;
  wire be_x_9_21;
  wire be_x_9_22;
  wire be_x_9_23;
  wire be_x_9_24;
  wire be_x_9_25;
  wire be_x_9_26;
  wire be_x_9_27;
  wire be_x_9_28;
  wire be_x_9_29;
  wire be_x_9_3;
  wire be_x_9_30;
  wire be_x_9_31;
  wire be_x_9_32;
  wire be_x_9_33;
  wire be_x_9_4;
  wire be_x_9_5;
  wire be_x_9_6;
  wire be_x_9_7;
  wire be_x_9_8;
  wire be_x_9_9;
  wire not_pp_0_35;
  wire not_pp_10_53;
  wire not_pp_11_55;
  wire not_pp_12_57;
  wire not_pp_13_59;
  wire not_pp_14_61;
  wire not_pp_15_63;
  wire not_pp_1_35;
  wire not_pp_2_37;
  wire not_pp_3_39;
  wire not_pp_4_41;
  wire not_pp_5_43;
  wire not_pp_6_45;
  wire not_pp_7_47;
  wire not_pp_8_49;
  wire not_pp_9_51;
  wire ny_0;
  wire ny_1;
  wire ny_10;
  wire ny_11;
  wire ny_12;
  wire ny_13;
  wire ny_14;
  wire ny_15;
  wire ny_16;
  wire ny_17;
  wire ny_18;
  wire ny_19;
  wire ny_2;
  wire ny_20;
  wire ny_21;
  wire ny_22;
  wire ny_23;
  wire ny_24;
  wire ny_25;
  wire ny_26;
  wire ny_27;
  wire ny_28;
  wire ny_29;
  wire ny_3;
  wire ny_30;
  wire ny_31;
  wire ny_4;
  wire ny_5;
  wire ny_6;
  wire ny_7;
  wire ny_8;
  wire ny_9;
  wire one;
  wire pp_0_0;
  wire pp_0_1;
  wire pp_0_10;
  wire pp_0_11;
  wire pp_0_12;
  wire pp_0_13;
  wire pp_0_14;
  wire pp_0_15;
  wire pp_0_16;
  wire pp_0_17;
  wire pp_0_18;
  wire pp_0_19;
  wire pp_0_2;
  wire pp_0_20;
  wire pp_0_21;
  wire pp_0_22;
  wire pp_0_23;
  wire pp_0_24;
  wire pp_0_25;
  wire pp_0_26;
  wire pp_0_27;
  wire pp_0_28;
  wire pp_0_29;
  wire pp_0_3;
  wire pp_0_30;
  wire pp_0_31;
  wire pp_0_32;
  wire pp_0_33;
  wire pp_0_4;
  wire pp_0_5;
  wire pp_0_6;
  wire pp_0_7;
  wire pp_0_8;
  wire pp_0_9;
  wire pp_10_20;
  wire pp_10_21;
  wire pp_10_22;
  wire pp_10_23;
  wire pp_10_24;
  wire pp_10_25;
  wire pp_10_26;
  wire pp_10_27;
  wire pp_10_28;
  wire pp_10_29;
  wire pp_10_30;
  wire pp_10_31;
  wire pp_10_32;
  wire pp_10_33;
  wire pp_10_34;
  wire pp_10_35;
  wire pp_10_36;
  wire pp_10_37;
  wire pp_10_38;
  wire pp_10_39;
  wire pp_10_40;
  wire pp_10_41;
  wire pp_10_42;
  wire pp_10_43;
  wire pp_10_44;
  wire pp_10_45;
  wire pp_10_46;
  wire pp_10_47;
  wire pp_10_48;
  wire pp_10_49;
  wire pp_10_50;
  wire pp_10_51;
  wire pp_10_52;
  wire pp_10_53;
  wire pp_11_22;
  wire pp_11_23;
  wire pp_11_24;
  wire pp_11_25;
  wire pp_11_26;
  wire pp_11_27;
  wire pp_11_28;
  wire pp_11_29;
  wire pp_11_30;
  wire pp_11_31;
  wire pp_11_32;
  wire pp_11_33;
  wire pp_11_34;
  wire pp_11_35;
  wire pp_11_36;
  wire pp_11_37;
  wire pp_11_38;
  wire pp_11_39;
  wire pp_11_40;
  wire pp_11_41;
  wire pp_11_42;
  wire pp_11_43;
  wire pp_11_44;
  wire pp_11_45;
  wire pp_11_46;
  wire pp_11_47;
  wire pp_11_48;
  wire pp_11_49;
  wire pp_11_50;
  wire pp_11_51;
  wire pp_11_52;
  wire pp_11_53;
  wire pp_11_54;
  wire pp_11_55;
  wire pp_12_24;
  wire pp_12_25;
  wire pp_12_26;
  wire pp_12_27;
  wire pp_12_28;
  wire pp_12_29;
  wire pp_12_30;
  wire pp_12_31;
  wire pp_12_32;
  wire pp_12_33;
  wire pp_12_34;
  wire pp_12_35;
  wire pp_12_36;
  wire pp_12_37;
  wire pp_12_38;
  wire pp_12_39;
  wire pp_12_40;
  wire pp_12_41;
  wire pp_12_42;
  wire pp_12_43;
  wire pp_12_44;
  wire pp_12_45;
  wire pp_12_46;
  wire pp_12_47;
  wire pp_12_48;
  wire pp_12_49;
  wire pp_12_50;
  wire pp_12_51;
  wire pp_12_52;
  wire pp_12_53;
  wire pp_12_54;
  wire pp_12_55;
  wire pp_12_56;
  wire pp_12_57;
  wire pp_13_26;
  wire pp_13_27;
  wire pp_13_28;
  wire pp_13_29;
  wire pp_13_30;
  wire pp_13_31;
  wire pp_13_32;
  wire pp_13_33;
  wire pp_13_34;
  wire pp_13_35;
  wire pp_13_36;
  wire pp_13_37;
  wire pp_13_38;
  wire pp_13_39;
  wire pp_13_40;
  wire pp_13_41;
  wire pp_13_42;
  wire pp_13_43;
  wire pp_13_44;
  wire pp_13_45;
  wire pp_13_46;
  wire pp_13_47;
  wire pp_13_48;
  wire pp_13_49;
  wire pp_13_50;
  wire pp_13_51;
  wire pp_13_52;
  wire pp_13_53;
  wire pp_13_54;
  wire pp_13_55;
  wire pp_13_56;
  wire pp_13_57;
  wire pp_13_58;
  wire pp_13_59;
  wire pp_14_28;
  wire pp_14_29;
  wire pp_14_30;
  wire pp_14_31;
  wire pp_14_32;
  wire pp_14_33;
  wire pp_14_34;
  wire pp_14_35;
  wire pp_14_36;
  wire pp_14_37;
  wire pp_14_38;
  wire pp_14_39;
  wire pp_14_40;
  wire pp_14_41;
  wire pp_14_42;
  wire pp_14_43;
  wire pp_14_44;
  wire pp_14_45;
  wire pp_14_46;
  wire pp_14_47;
  wire pp_14_48;
  wire pp_14_49;
  wire pp_14_50;
  wire pp_14_51;
  wire pp_14_52;
  wire pp_14_53;
  wire pp_14_54;
  wire pp_14_55;
  wire pp_14_56;
  wire pp_14_57;
  wire pp_14_58;
  wire pp_14_59;
  wire pp_14_60;
  wire pp_14_61;
  wire pp_15_30;
  wire pp_15_31;
  wire pp_15_32;
  wire pp_15_33;
  wire pp_15_34;
  wire pp_15_35;
  wire pp_15_36;
  wire pp_15_37;
  wire pp_15_38;
  wire pp_15_39;
  wire pp_15_40;
  wire pp_15_41;
  wire pp_15_42;
  wire pp_15_43;
  wire pp_15_44;
  wire pp_15_45;
  wire pp_15_46;
  wire pp_15_47;
  wire pp_15_48;
  wire pp_15_49;
  wire pp_15_50;
  wire pp_15_51;
  wire pp_15_52;
  wire pp_15_53;
  wire pp_15_54;
  wire pp_15_55;
  wire pp_15_56;
  wire pp_15_57;
  wire pp_15_58;
  wire pp_15_59;
  wire pp_15_60;
  wire pp_15_61;
  wire pp_15_62;
  wire pp_15_63;
  wire pp_16_32;
  wire pp_16_33;
  wire pp_16_34;
  wire pp_16_35;
  wire pp_16_36;
  wire pp_16_37;
  wire pp_16_38;
  wire pp_16_39;
  wire pp_16_40;
  wire pp_16_41;
  wire pp_16_42;
  wire pp_16_43;
  wire pp_16_44;
  wire pp_16_45;
  wire pp_16_46;
  wire pp_16_47;
  wire pp_16_48;
  wire pp_16_49;
  wire pp_16_50;
  wire pp_16_51;
  wire pp_16_52;
  wire pp_16_53;
  wire pp_16_54;
  wire pp_16_55;
  wire pp_16_56;
  wire pp_16_57;
  wire pp_16_58;
  wire pp_16_59;
  wire pp_16_60;
  wire pp_16_61;
  wire pp_16_62;
  wire pp_16_63;
  wire pp_1_10;
  wire pp_1_11;
  wire pp_1_12;
  wire pp_1_13;
  wire pp_1_14;
  wire pp_1_15;
  wire pp_1_16;
  wire pp_1_17;
  wire pp_1_18;
  wire pp_1_19;
  wire pp_1_2;
  wire pp_1_20;
  wire pp_1_21;
  wire pp_1_22;
  wire pp_1_23;
  wire pp_1_24;
  wire pp_1_25;
  wire pp_1_26;
  wire pp_1_27;
  wire pp_1_28;
  wire pp_1_29;
  wire pp_1_3;
  wire pp_1_30;
  wire pp_1_31;
  wire pp_1_32;
  wire pp_1_33;
  wire pp_1_34;
  wire pp_1_35;
  wire pp_1_4;
  wire pp_1_5;
  wire pp_1_6;
  wire pp_1_7;
  wire pp_1_8;
  wire pp_1_9;
  wire pp_2_10;
  wire pp_2_11;
  wire pp_2_12;
  wire pp_2_13;
  wire pp_2_14;
  wire pp_2_15;
  wire pp_2_16;
  wire pp_2_17;
  wire pp_2_18;
  wire pp_2_19;
  wire pp_2_20;
  wire pp_2_21;
  wire pp_2_22;
  wire pp_2_23;
  wire pp_2_24;
  wire pp_2_25;
  wire pp_2_26;
  wire pp_2_27;
  wire pp_2_28;
  wire pp_2_29;
  wire pp_2_30;
  wire pp_2_31;
  wire pp_2_32;
  wire pp_2_33;
  wire pp_2_34;
  wire pp_2_35;
  wire pp_2_36;
  wire pp_2_37;
  wire pp_2_4;
  wire pp_2_5;
  wire pp_2_6;
  wire pp_2_7;
  wire pp_2_8;
  wire pp_2_9;
  wire pp_3_10;
  wire pp_3_11;
  wire pp_3_12;
  wire pp_3_13;
  wire pp_3_14;
  wire pp_3_15;
  wire pp_3_16;
  wire pp_3_17;
  wire pp_3_18;
  wire pp_3_19;
  wire pp_3_20;
  wire pp_3_21;
  wire pp_3_22;
  wire pp_3_23;
  wire pp_3_24;
  wire pp_3_25;
  wire pp_3_26;
  wire pp_3_27;
  wire pp_3_28;
  wire pp_3_29;
  wire pp_3_30;
  wire pp_3_31;
  wire pp_3_32;
  wire pp_3_33;
  wire pp_3_34;
  wire pp_3_35;
  wire pp_3_36;
  wire pp_3_37;
  wire pp_3_38;
  wire pp_3_39;
  wire pp_3_6;
  wire pp_3_7;
  wire pp_3_8;
  wire pp_3_9;
  wire pp_4_10;
  wire pp_4_11;
  wire pp_4_12;
  wire pp_4_13;
  wire pp_4_14;
  wire pp_4_15;
  wire pp_4_16;
  wire pp_4_17;
  wire pp_4_18;
  wire pp_4_19;
  wire pp_4_20;
  wire pp_4_21;
  wire pp_4_22;
  wire pp_4_23;
  wire pp_4_24;
  wire pp_4_25;
  wire pp_4_26;
  wire pp_4_27;
  wire pp_4_28;
  wire pp_4_29;
  wire pp_4_30;
  wire pp_4_31;
  wire pp_4_32;
  wire pp_4_33;
  wire pp_4_34;
  wire pp_4_35;
  wire pp_4_36;
  wire pp_4_37;
  wire pp_4_38;
  wire pp_4_39;
  wire pp_4_40;
  wire pp_4_41;
  wire pp_4_8;
  wire pp_4_9;
  wire pp_5_10;
  wire pp_5_11;
  wire pp_5_12;
  wire pp_5_13;
  wire pp_5_14;
  wire pp_5_15;
  wire pp_5_16;
  wire pp_5_17;
  wire pp_5_18;
  wire pp_5_19;
  wire pp_5_20;
  wire pp_5_21;
  wire pp_5_22;
  wire pp_5_23;
  wire pp_5_24;
  wire pp_5_25;
  wire pp_5_26;
  wire pp_5_27;
  wire pp_5_28;
  wire pp_5_29;
  wire pp_5_30;
  wire pp_5_31;
  wire pp_5_32;
  wire pp_5_33;
  wire pp_5_34;
  wire pp_5_35;
  wire pp_5_36;
  wire pp_5_37;
  wire pp_5_38;
  wire pp_5_39;
  wire pp_5_40;
  wire pp_5_41;
  wire pp_5_42;
  wire pp_5_43;
  wire pp_6_12;
  wire pp_6_13;
  wire pp_6_14;
  wire pp_6_15;
  wire pp_6_16;
  wire pp_6_17;
  wire pp_6_18;
  wire pp_6_19;
  wire pp_6_20;
  wire pp_6_21;
  wire pp_6_22;
  wire pp_6_23;
  wire pp_6_24;
  wire pp_6_25;
  wire pp_6_26;
  wire pp_6_27;
  wire pp_6_28;
  wire pp_6_29;
  wire pp_6_30;
  wire pp_6_31;
  wire pp_6_32;
  wire pp_6_33;
  wire pp_6_34;
  wire pp_6_35;
  wire pp_6_36;
  wire pp_6_37;
  wire pp_6_38;
  wire pp_6_39;
  wire pp_6_40;
  wire pp_6_41;
  wire pp_6_42;
  wire pp_6_43;
  wire pp_6_44;
  wire pp_6_45;
  wire pp_7_14;
  wire pp_7_15;
  wire pp_7_16;
  wire pp_7_17;
  wire pp_7_18;
  wire pp_7_19;
  wire pp_7_20;
  wire pp_7_21;
  wire pp_7_22;
  wire pp_7_23;
  wire pp_7_24;
  wire pp_7_25;
  wire pp_7_26;
  wire pp_7_27;
  wire pp_7_28;
  wire pp_7_29;
  wire pp_7_30;
  wire pp_7_31;
  wire pp_7_32;
  wire pp_7_33;
  wire pp_7_34;
  wire pp_7_35;
  wire pp_7_36;
  wire pp_7_37;
  wire pp_7_38;
  wire pp_7_39;
  wire pp_7_40;
  wire pp_7_41;
  wire pp_7_42;
  wire pp_7_43;
  wire pp_7_44;
  wire pp_7_45;
  wire pp_7_46;
  wire pp_7_47;
  wire pp_8_16;
  wire pp_8_17;
  wire pp_8_18;
  wire pp_8_19;
  wire pp_8_20;
  wire pp_8_21;
  wire pp_8_22;
  wire pp_8_23;
  wire pp_8_24;
  wire pp_8_25;
  wire pp_8_26;
  wire pp_8_27;
  wire pp_8_28;
  wire pp_8_29;
  wire pp_8_30;
  wire pp_8_31;
  wire pp_8_32;
  wire pp_8_33;
  wire pp_8_34;
  wire pp_8_35;
  wire pp_8_36;
  wire pp_8_37;
  wire pp_8_38;
  wire pp_8_39;
  wire pp_8_40;
  wire pp_8_41;
  wire pp_8_42;
  wire pp_8_43;
  wire pp_8_44;
  wire pp_8_45;
  wire pp_8_46;
  wire pp_8_47;
  wire pp_8_48;
  wire pp_8_49;
  wire pp_9_18;
  wire pp_9_19;
  wire pp_9_20;
  wire pp_9_21;
  wire pp_9_22;
  wire pp_9_23;
  wire pp_9_24;
  wire pp_9_25;
  wire pp_9_26;
  wire pp_9_27;
  wire pp_9_28;
  wire pp_9_29;
  wire pp_9_30;
  wire pp_9_31;
  wire pp_9_32;
  wire pp_9_33;
  wire pp_9_34;
  wire pp_9_35;
  wire pp_9_36;
  wire pp_9_37;
  wire pp_9_38;
  wire pp_9_39;
  wire pp_9_40;
  wire pp_9_41;
  wire pp_9_42;
  wire pp_9_43;
  wire pp_9_44;
  wire pp_9_45;
  wire pp_9_46;
  wire pp_9_47;
  wire pp_9_48;
  wire pp_9_49;
  wire pp_9_50;
  wire pp_9_51;
  wire px_0_0;
  wire px_0_1;
  wire px_0_10;
  wire px_0_11;
  wire px_0_12;
  wire px_0_13;
  wire px_0_14;
  wire px_0_15;
  wire px_0_16;
  wire px_0_17;
  wire px_0_18;
  wire px_0_19;
  wire px_0_2;
  wire px_0_20;
  wire px_0_21;
  wire px_0_22;
  wire px_0_23;
  wire px_0_24;
  wire px_0_25;
  wire px_0_26;
  wire px_0_27;
  wire px_0_28;
  wire px_0_29;
  wire px_0_3;
  wire px_0_30;
  wire px_0_31;
  wire px_0_32;
  wire px_0_33;
  wire px_0_34;
  wire px_0_4;
  wire px_0_5;
  wire px_0_6;
  wire px_0_7;
  wire px_0_8;
  wire px_0_9;
  wire px_10_0;
  wire px_10_1;
  wire px_10_10;
  wire px_10_11;
  wire px_10_12;
  wire px_10_13;
  wire px_10_14;
  wire px_10_15;
  wire px_10_16;
  wire px_10_17;
  wire px_10_18;
  wire px_10_19;
  wire px_10_2;
  wire px_10_20;
  wire px_10_21;
  wire px_10_22;
  wire px_10_23;
  wire px_10_24;
  wire px_10_25;
  wire px_10_26;
  wire px_10_27;
  wire px_10_28;
  wire px_10_29;
  wire px_10_3;
  wire px_10_30;
  wire px_10_31;
  wire px_10_32;
  wire px_10_33;
  wire px_10_34;
  wire px_10_4;
  wire px_10_5;
  wire px_10_6;
  wire px_10_7;
  wire px_10_8;
  wire px_10_9;
  wire px_11_0;
  wire px_11_1;
  wire px_11_10;
  wire px_11_11;
  wire px_11_12;
  wire px_11_13;
  wire px_11_14;
  wire px_11_15;
  wire px_11_16;
  wire px_11_17;
  wire px_11_18;
  wire px_11_19;
  wire px_11_2;
  wire px_11_20;
  wire px_11_21;
  wire px_11_22;
  wire px_11_23;
  wire px_11_24;
  wire px_11_25;
  wire px_11_26;
  wire px_11_27;
  wire px_11_28;
  wire px_11_29;
  wire px_11_3;
  wire px_11_30;
  wire px_11_31;
  wire px_11_32;
  wire px_11_33;
  wire px_11_34;
  wire px_11_4;
  wire px_11_5;
  wire px_11_6;
  wire px_11_7;
  wire px_11_8;
  wire px_11_9;
  wire px_12_0;
  wire px_12_1;
  wire px_12_10;
  wire px_12_11;
  wire px_12_12;
  wire px_12_13;
  wire px_12_14;
  wire px_12_15;
  wire px_12_16;
  wire px_12_17;
  wire px_12_18;
  wire px_12_19;
  wire px_12_2;
  wire px_12_20;
  wire px_12_21;
  wire px_12_22;
  wire px_12_23;
  wire px_12_24;
  wire px_12_25;
  wire px_12_26;
  wire px_12_27;
  wire px_12_28;
  wire px_12_29;
  wire px_12_3;
  wire px_12_30;
  wire px_12_31;
  wire px_12_32;
  wire px_12_33;
  wire px_12_34;
  wire px_12_4;
  wire px_12_5;
  wire px_12_6;
  wire px_12_7;
  wire px_12_8;
  wire px_12_9;
  wire px_13_0;
  wire px_13_1;
  wire px_13_10;
  wire px_13_11;
  wire px_13_12;
  wire px_13_13;
  wire px_13_14;
  wire px_13_15;
  wire px_13_16;
  wire px_13_17;
  wire px_13_18;
  wire px_13_19;
  wire px_13_2;
  wire px_13_20;
  wire px_13_21;
  wire px_13_22;
  wire px_13_23;
  wire px_13_24;
  wire px_13_25;
  wire px_13_26;
  wire px_13_27;
  wire px_13_28;
  wire px_13_29;
  wire px_13_3;
  wire px_13_30;
  wire px_13_31;
  wire px_13_32;
  wire px_13_33;
  wire px_13_34;
  wire px_13_4;
  wire px_13_5;
  wire px_13_6;
  wire px_13_7;
  wire px_13_8;
  wire px_13_9;
  wire px_14_0;
  wire px_14_1;
  wire px_14_10;
  wire px_14_11;
  wire px_14_12;
  wire px_14_13;
  wire px_14_14;
  wire px_14_15;
  wire px_14_16;
  wire px_14_17;
  wire px_14_18;
  wire px_14_19;
  wire px_14_2;
  wire px_14_20;
  wire px_14_21;
  wire px_14_22;
  wire px_14_23;
  wire px_14_24;
  wire px_14_25;
  wire px_14_26;
  wire px_14_27;
  wire px_14_28;
  wire px_14_29;
  wire px_14_3;
  wire px_14_30;
  wire px_14_31;
  wire px_14_32;
  wire px_14_33;
  wire px_14_34;
  wire px_14_4;
  wire px_14_5;
  wire px_14_6;
  wire px_14_7;
  wire px_14_8;
  wire px_14_9;
  wire px_15_0;
  wire px_15_1;
  wire px_15_10;
  wire px_15_11;
  wire px_15_12;
  wire px_15_13;
  wire px_15_14;
  wire px_15_15;
  wire px_15_16;
  wire px_15_17;
  wire px_15_18;
  wire px_15_19;
  wire px_15_2;
  wire px_15_20;
  wire px_15_21;
  wire px_15_22;
  wire px_15_23;
  wire px_15_24;
  wire px_15_25;
  wire px_15_26;
  wire px_15_27;
  wire px_15_28;
  wire px_15_29;
  wire px_15_3;
  wire px_15_30;
  wire px_15_31;
  wire px_15_32;
  wire px_15_33;
  wire px_15_34;
  wire px_15_4;
  wire px_15_5;
  wire px_15_6;
  wire px_15_7;
  wire px_15_8;
  wire px_15_9;
  wire px_16_0;
  wire px_16_1;
  wire px_16_10;
  wire px_16_11;
  wire px_16_12;
  wire px_16_13;
  wire px_16_14;
  wire px_16_15;
  wire px_16_16;
  wire px_16_17;
  wire px_16_18;
  wire px_16_19;
  wire px_16_2;
  wire px_16_20;
  wire px_16_21;
  wire px_16_22;
  wire px_16_23;
  wire px_16_24;
  wire px_16_25;
  wire px_16_26;
  wire px_16_27;
  wire px_16_28;
  wire px_16_29;
  wire px_16_3;
  wire px_16_30;
  wire px_16_31;
  wire px_16_32;
  wire px_16_33;
  wire px_16_34;
  wire px_16_4;
  wire px_16_5;
  wire px_16_6;
  wire px_16_7;
  wire px_16_8;
  wire px_16_9;
  wire px_1_0;
  wire px_1_1;
  wire px_1_10;
  wire px_1_11;
  wire px_1_12;
  wire px_1_13;
  wire px_1_14;
  wire px_1_15;
  wire px_1_16;
  wire px_1_17;
  wire px_1_18;
  wire px_1_19;
  wire px_1_2;
  wire px_1_20;
  wire px_1_21;
  wire px_1_22;
  wire px_1_23;
  wire px_1_24;
  wire px_1_25;
  wire px_1_26;
  wire px_1_27;
  wire px_1_28;
  wire px_1_29;
  wire px_1_3;
  wire px_1_30;
  wire px_1_31;
  wire px_1_32;
  wire px_1_33;
  wire px_1_34;
  wire px_1_4;
  wire px_1_5;
  wire px_1_6;
  wire px_1_7;
  wire px_1_8;
  wire px_1_9;
  wire px_2_0;
  wire px_2_1;
  wire px_2_10;
  wire px_2_11;
  wire px_2_12;
  wire px_2_13;
  wire px_2_14;
  wire px_2_15;
  wire px_2_16;
  wire px_2_17;
  wire px_2_18;
  wire px_2_19;
  wire px_2_2;
  wire px_2_20;
  wire px_2_21;
  wire px_2_22;
  wire px_2_23;
  wire px_2_24;
  wire px_2_25;
  wire px_2_26;
  wire px_2_27;
  wire px_2_28;
  wire px_2_29;
  wire px_2_3;
  wire px_2_30;
  wire px_2_31;
  wire px_2_32;
  wire px_2_33;
  wire px_2_34;
  wire px_2_4;
  wire px_2_5;
  wire px_2_6;
  wire px_2_7;
  wire px_2_8;
  wire px_2_9;
  wire px_3_0;
  wire px_3_1;
  wire px_3_10;
  wire px_3_11;
  wire px_3_12;
  wire px_3_13;
  wire px_3_14;
  wire px_3_15;
  wire px_3_16;
  wire px_3_17;
  wire px_3_18;
  wire px_3_19;
  wire px_3_2;
  wire px_3_20;
  wire px_3_21;
  wire px_3_22;
  wire px_3_23;
  wire px_3_24;
  wire px_3_25;
  wire px_3_26;
  wire px_3_27;
  wire px_3_28;
  wire px_3_29;
  wire px_3_3;
  wire px_3_30;
  wire px_3_31;
  wire px_3_32;
  wire px_3_33;
  wire px_3_34;
  wire px_3_4;
  wire px_3_5;
  wire px_3_6;
  wire px_3_7;
  wire px_3_8;
  wire px_3_9;
  wire px_4_0;
  wire px_4_1;
  wire px_4_10;
  wire px_4_11;
  wire px_4_12;
  wire px_4_13;
  wire px_4_14;
  wire px_4_15;
  wire px_4_16;
  wire px_4_17;
  wire px_4_18;
  wire px_4_19;
  wire px_4_2;
  wire px_4_20;
  wire px_4_21;
  wire px_4_22;
  wire px_4_23;
  wire px_4_24;
  wire px_4_25;
  wire px_4_26;
  wire px_4_27;
  wire px_4_28;
  wire px_4_29;
  wire px_4_3;
  wire px_4_30;
  wire px_4_31;
  wire px_4_32;
  wire px_4_33;
  wire px_4_34;
  wire px_4_4;
  wire px_4_5;
  wire px_4_6;
  wire px_4_7;
  wire px_4_8;
  wire px_4_9;
  wire px_5_0;
  wire px_5_1;
  wire px_5_10;
  wire px_5_11;
  wire px_5_12;
  wire px_5_13;
  wire px_5_14;
  wire px_5_15;
  wire px_5_16;
  wire px_5_17;
  wire px_5_18;
  wire px_5_19;
  wire px_5_2;
  wire px_5_20;
  wire px_5_21;
  wire px_5_22;
  wire px_5_23;
  wire px_5_24;
  wire px_5_25;
  wire px_5_26;
  wire px_5_27;
  wire px_5_28;
  wire px_5_29;
  wire px_5_3;
  wire px_5_30;
  wire px_5_31;
  wire px_5_32;
  wire px_5_33;
  wire px_5_34;
  wire px_5_4;
  wire px_5_5;
  wire px_5_6;
  wire px_5_7;
  wire px_5_8;
  wire px_5_9;
  wire px_6_0;
  wire px_6_1;
  wire px_6_10;
  wire px_6_11;
  wire px_6_12;
  wire px_6_13;
  wire px_6_14;
  wire px_6_15;
  wire px_6_16;
  wire px_6_17;
  wire px_6_18;
  wire px_6_19;
  wire px_6_2;
  wire px_6_20;
  wire px_6_21;
  wire px_6_22;
  wire px_6_23;
  wire px_6_24;
  wire px_6_25;
  wire px_6_26;
  wire px_6_27;
  wire px_6_28;
  wire px_6_29;
  wire px_6_3;
  wire px_6_30;
  wire px_6_31;
  wire px_6_32;
  wire px_6_33;
  wire px_6_34;
  wire px_6_4;
  wire px_6_5;
  wire px_6_6;
  wire px_6_7;
  wire px_6_8;
  wire px_6_9;
  wire px_7_0;
  wire px_7_1;
  wire px_7_10;
  wire px_7_11;
  wire px_7_12;
  wire px_7_13;
  wire px_7_14;
  wire px_7_15;
  wire px_7_16;
  wire px_7_17;
  wire px_7_18;
  wire px_7_19;
  wire px_7_2;
  wire px_7_20;
  wire px_7_21;
  wire px_7_22;
  wire px_7_23;
  wire px_7_24;
  wire px_7_25;
  wire px_7_26;
  wire px_7_27;
  wire px_7_28;
  wire px_7_29;
  wire px_7_3;
  wire px_7_30;
  wire px_7_31;
  wire px_7_32;
  wire px_7_33;
  wire px_7_34;
  wire px_7_4;
  wire px_7_5;
  wire px_7_6;
  wire px_7_7;
  wire px_7_8;
  wire px_7_9;
  wire px_8_0;
  wire px_8_1;
  wire px_8_10;
  wire px_8_11;
  wire px_8_12;
  wire px_8_13;
  wire px_8_14;
  wire px_8_15;
  wire px_8_16;
  wire px_8_17;
  wire px_8_18;
  wire px_8_19;
  wire px_8_2;
  wire px_8_20;
  wire px_8_21;
  wire px_8_22;
  wire px_8_23;
  wire px_8_24;
  wire px_8_25;
  wire px_8_26;
  wire px_8_27;
  wire px_8_28;
  wire px_8_29;
  wire px_8_3;
  wire px_8_30;
  wire px_8_31;
  wire px_8_32;
  wire px_8_33;
  wire px_8_34;
  wire px_8_4;
  wire px_8_5;
  wire px_8_6;
  wire px_8_7;
  wire px_8_8;
  wire px_8_9;
  wire px_9_0;
  wire px_9_1;
  wire px_9_10;
  wire px_9_11;
  wire px_9_12;
  wire px_9_13;
  wire px_9_14;
  wire px_9_15;
  wire px_9_16;
  wire px_9_17;
  wire px_9_18;
  wire px_9_19;
  wire px_9_2;
  wire px_9_20;
  wire px_9_21;
  wire px_9_22;
  wire px_9_23;
  wire px_9_24;
  wire px_9_25;
  wire px_9_26;
  wire px_9_27;
  wire px_9_28;
  wire px_9_29;
  wire px_9_3;
  wire px_9_30;
  wire px_9_31;
  wire px_9_32;
  wire px_9_33;
  wire px_9_34;
  wire px_9_4;
  wire px_9_5;
  wire px_9_6;
  wire px_9_7;
  wire px_9_8;
  wire px_9_9;
  wire x_0;
  wire x_1;
  wire x_10;
  wire x_11;
  wire x_12;
  wire x_13;
  wire x_14;
  wire x_15;
  wire x_16;
  wire x_17;
  wire x_18;
  wire x_19;
  wire x_2;
  wire x_20;
  wire x_21;
  wire x_22;
  wire x_23;
  wire x_24;
  wire x_25;
  wire x_26;
  wire x_27;
  wire x_28;
  wire x_29;
  wire x_3;
  wire x_30;
  wire x_31;
  wire x_4;
  wire x_5;
  wire x_6;
  wire x_7;
  wire x_8;
  wire x_9;
  wire y_0;
  wire y_1;
  wire y_10;
  wire y_11;
  wire y_12;
  wire y_13;
  wire y_14;
  wire y_15;
  wire y_16;
  wire y_17;
  wire y_18;
  wire y_19;
  wire y_2;
  wire y_20;
  wire y_21;
  wire y_22;
  wire y_23;
  wire y_24;
  wire y_25;
  wire y_26;
  wire y_27;
  wire y_28;
  wire y_29;
  wire y_3;
  wire y_30;
  wire y_31;
  wire y_4;
  wire y_5;
  wire y_6;
  wire y_7;
  wire y_8;
  wire y_9;
  wire zero;
  assign be_2x_0_0 = ~(px_0_0 & be_s2_0);
  assign be_2x_0_1 = ~(px_0_1 & be_s2_0);
  assign be_2x_0_10 = ~(px_0_10 & be_s2_0);
  assign be_2x_0_11 = ~(px_0_11 & be_s2_0);
  assign be_2x_0_12 = ~(px_0_12 & be_s2_0);
  assign be_2x_0_13 = ~(px_0_13 & be_s2_0);
  assign be_2x_0_14 = ~(px_0_14 & be_s2_0);
  assign be_2x_0_15 = ~(px_0_15 & be_s2_0);
  assign be_2x_0_16 = ~(px_0_16 & be_s2_0);
  assign be_2x_0_17 = ~(px_0_17 & be_s2_0);
  assign be_2x_0_18 = ~(px_0_18 & be_s2_0);
  assign be_2x_0_19 = ~(px_0_19 & be_s2_0);
  assign be_2x_0_2 = ~(px_0_2 & be_s2_0);
  assign be_2x_0_20 = ~(px_0_20 & be_s2_0);
  assign be_2x_0_21 = ~(px_0_21 & be_s2_0);
  assign be_2x_0_22 = ~(px_0_22 & be_s2_0);
  assign be_2x_0_23 = ~(px_0_23 & be_s2_0);
  assign be_2x_0_24 = ~(px_0_24 & be_s2_0);
  assign be_2x_0_25 = ~(px_0_25 & be_s2_0);
  assign be_2x_0_26 = ~(px_0_26 & be_s2_0);
  assign be_2x_0_27 = ~(px_0_27 & be_s2_0);
  assign be_2x_0_28 = ~(px_0_28 & be_s2_0);
  assign be_2x_0_29 = ~(px_0_29 & be_s2_0);
  assign be_2x_0_3 = ~(px_0_3 & be_s2_0);
  assign be_2x_0_30 = ~(px_0_30 & be_s2_0);
  assign be_2x_0_31 = ~(px_0_31 & be_s2_0);
  assign be_2x_0_32 = ~(px_0_32 & be_s2_0);
  assign be_2x_0_33 = ~(px_0_33 & be_s2_0);
  assign be_2x_0_4 = ~(px_0_4 & be_s2_0);
  assign be_2x_0_5 = ~(px_0_5 & be_s2_0);
  assign be_2x_0_6 = ~(px_0_6 & be_s2_0);
  assign be_2x_0_7 = ~(px_0_7 & be_s2_0);
  assign be_2x_0_8 = ~(px_0_8 & be_s2_0);
  assign be_2x_0_9 = ~(px_0_9 & be_s2_0);
  assign be_2x_10_0 = ~(px_10_0 & be_s2_10);
  assign be_2x_10_1 = ~(px_10_1 & be_s2_10);
  assign be_2x_10_10 = ~(px_10_10 & be_s2_10);
  assign be_2x_10_11 = ~(px_10_11 & be_s2_10);
  assign be_2x_10_12 = ~(px_10_12 & be_s2_10);
  assign be_2x_10_13 = ~(px_10_13 & be_s2_10);
  assign be_2x_10_14 = ~(px_10_14 & be_s2_10);
  assign be_2x_10_15 = ~(px_10_15 & be_s2_10);
  assign be_2x_10_16 = ~(px_10_16 & be_s2_10);
  assign be_2x_10_17 = ~(px_10_17 & be_s2_10);
  assign be_2x_10_18 = ~(px_10_18 & be_s2_10);
  assign be_2x_10_19 = ~(px_10_19 & be_s2_10);
  assign be_2x_10_2 = ~(px_10_2 & be_s2_10);
  assign be_2x_10_20 = ~(px_10_20 & be_s2_10);
  assign be_2x_10_21 = ~(px_10_21 & be_s2_10);
  assign be_2x_10_22 = ~(px_10_22 & be_s2_10);
  assign be_2x_10_23 = ~(px_10_23 & be_s2_10);
  assign be_2x_10_24 = ~(px_10_24 & be_s2_10);
  assign be_2x_10_25 = ~(px_10_25 & be_s2_10);
  assign be_2x_10_26 = ~(px_10_26 & be_s2_10);
  assign be_2x_10_27 = ~(px_10_27 & be_s2_10);
  assign be_2x_10_28 = ~(px_10_28 & be_s2_10);
  assign be_2x_10_29 = ~(px_10_29 & be_s2_10);
  assign be_2x_10_3 = ~(px_10_3 & be_s2_10);
  assign be_2x_10_30 = ~(px_10_30 & be_s2_10);
  assign be_2x_10_31 = ~(px_10_31 & be_s2_10);
  assign be_2x_10_32 = ~(px_10_32 & be_s2_10);
  assign be_2x_10_33 = ~(px_10_33 & be_s2_10);
  assign be_2x_10_4 = ~(px_10_4 & be_s2_10);
  assign be_2x_10_5 = ~(px_10_5 & be_s2_10);
  assign be_2x_10_6 = ~(px_10_6 & be_s2_10);
  assign be_2x_10_7 = ~(px_10_7 & be_s2_10);
  assign be_2x_10_8 = ~(px_10_8 & be_s2_10);
  assign be_2x_10_9 = ~(px_10_9 & be_s2_10);
  assign be_2x_11_0 = ~(px_11_0 & be_s2_11);
  assign be_2x_11_1 = ~(px_11_1 & be_s2_11);
  assign be_2x_11_10 = ~(px_11_10 & be_s2_11);
  assign be_2x_11_11 = ~(px_11_11 & be_s2_11);
  assign be_2x_11_12 = ~(px_11_12 & be_s2_11);
  assign be_2x_11_13 = ~(px_11_13 & be_s2_11);
  assign be_2x_11_14 = ~(px_11_14 & be_s2_11);
  assign be_2x_11_15 = ~(px_11_15 & be_s2_11);
  assign be_2x_11_16 = ~(px_11_16 & be_s2_11);
  assign be_2x_11_17 = ~(px_11_17 & be_s2_11);
  assign be_2x_11_18 = ~(px_11_18 & be_s2_11);
  assign be_2x_11_19 = ~(px_11_19 & be_s2_11);
  assign be_2x_11_2 = ~(px_11_2 & be_s2_11);
  assign be_2x_11_20 = ~(px_11_20 & be_s2_11);
  assign be_2x_11_21 = ~(px_11_21 & be_s2_11);
  assign be_2x_11_22 = ~(px_11_22 & be_s2_11);
  assign be_2x_11_23 = ~(px_11_23 & be_s2_11);
  assign be_2x_11_24 = ~(px_11_24 & be_s2_11);
  assign be_2x_11_25 = ~(px_11_25 & be_s2_11);
  assign be_2x_11_26 = ~(px_11_26 & be_s2_11);
  assign be_2x_11_27 = ~(px_11_27 & be_s2_11);
  assign be_2x_11_28 = ~(px_11_28 & be_s2_11);
  assign be_2x_11_29 = ~(px_11_29 & be_s2_11);
  assign be_2x_11_3 = ~(px_11_3 & be_s2_11);
  assign be_2x_11_30 = ~(px_11_30 & be_s2_11);
  assign be_2x_11_31 = ~(px_11_31 & be_s2_11);
  assign be_2x_11_32 = ~(px_11_32 & be_s2_11);
  assign be_2x_11_33 = ~(px_11_33 & be_s2_11);
  assign be_2x_11_4 = ~(px_11_4 & be_s2_11);
  assign be_2x_11_5 = ~(px_11_5 & be_s2_11);
  assign be_2x_11_6 = ~(px_11_6 & be_s2_11);
  assign be_2x_11_7 = ~(px_11_7 & be_s2_11);
  assign be_2x_11_8 = ~(px_11_8 & be_s2_11);
  assign be_2x_11_9 = ~(px_11_9 & be_s2_11);
  assign be_2x_12_0 = ~(px_12_0 & be_s2_12);
  assign be_2x_12_1 = ~(px_12_1 & be_s2_12);
  assign be_2x_12_10 = ~(px_12_10 & be_s2_12);
  assign be_2x_12_11 = ~(px_12_11 & be_s2_12);
  assign be_2x_12_12 = ~(px_12_12 & be_s2_12);
  assign be_2x_12_13 = ~(px_12_13 & be_s2_12);
  assign be_2x_12_14 = ~(px_12_14 & be_s2_12);
  assign be_2x_12_15 = ~(px_12_15 & be_s2_12);
  assign be_2x_12_16 = ~(px_12_16 & be_s2_12);
  assign be_2x_12_17 = ~(px_12_17 & be_s2_12);
  assign be_2x_12_18 = ~(px_12_18 & be_s2_12);
  assign be_2x_12_19 = ~(px_12_19 & be_s2_12);
  assign be_2x_12_2 = ~(px_12_2 & be_s2_12);
  assign be_2x_12_20 = ~(px_12_20 & be_s2_12);
  assign be_2x_12_21 = ~(px_12_21 & be_s2_12);
  assign be_2x_12_22 = ~(px_12_22 & be_s2_12);
  assign be_2x_12_23 = ~(px_12_23 & be_s2_12);
  assign be_2x_12_24 = ~(px_12_24 & be_s2_12);
  assign be_2x_12_25 = ~(px_12_25 & be_s2_12);
  assign be_2x_12_26 = ~(px_12_26 & be_s2_12);
  assign be_2x_12_27 = ~(px_12_27 & be_s2_12);
  assign be_2x_12_28 = ~(px_12_28 & be_s2_12);
  assign be_2x_12_29 = ~(px_12_29 & be_s2_12);
  assign be_2x_12_3 = ~(px_12_3 & be_s2_12);
  assign be_2x_12_30 = ~(px_12_30 & be_s2_12);
  assign be_2x_12_31 = ~(px_12_31 & be_s2_12);
  assign be_2x_12_32 = ~(px_12_32 & be_s2_12);
  assign be_2x_12_33 = ~(px_12_33 & be_s2_12);
  assign be_2x_12_4 = ~(px_12_4 & be_s2_12);
  assign be_2x_12_5 = ~(px_12_5 & be_s2_12);
  assign be_2x_12_6 = ~(px_12_6 & be_s2_12);
  assign be_2x_12_7 = ~(px_12_7 & be_s2_12);
  assign be_2x_12_8 = ~(px_12_8 & be_s2_12);
  assign be_2x_12_9 = ~(px_12_9 & be_s2_12);
  assign be_2x_13_0 = ~(px_13_0 & be_s2_13);
  assign be_2x_13_1 = ~(px_13_1 & be_s2_13);
  assign be_2x_13_10 = ~(px_13_10 & be_s2_13);
  assign be_2x_13_11 = ~(px_13_11 & be_s2_13);
  assign be_2x_13_12 = ~(px_13_12 & be_s2_13);
  assign be_2x_13_13 = ~(px_13_13 & be_s2_13);
  assign be_2x_13_14 = ~(px_13_14 & be_s2_13);
  assign be_2x_13_15 = ~(px_13_15 & be_s2_13);
  assign be_2x_13_16 = ~(px_13_16 & be_s2_13);
  assign be_2x_13_17 = ~(px_13_17 & be_s2_13);
  assign be_2x_13_18 = ~(px_13_18 & be_s2_13);
  assign be_2x_13_19 = ~(px_13_19 & be_s2_13);
  assign be_2x_13_2 = ~(px_13_2 & be_s2_13);
  assign be_2x_13_20 = ~(px_13_20 & be_s2_13);
  assign be_2x_13_21 = ~(px_13_21 & be_s2_13);
  assign be_2x_13_22 = ~(px_13_22 & be_s2_13);
  assign be_2x_13_23 = ~(px_13_23 & be_s2_13);
  assign be_2x_13_24 = ~(px_13_24 & be_s2_13);
  assign be_2x_13_25 = ~(px_13_25 & be_s2_13);
  assign be_2x_13_26 = ~(px_13_26 & be_s2_13);
  assign be_2x_13_27 = ~(px_13_27 & be_s2_13);
  assign be_2x_13_28 = ~(px_13_28 & be_s2_13);
  assign be_2x_13_29 = ~(px_13_29 & be_s2_13);
  assign be_2x_13_3 = ~(px_13_3 & be_s2_13);
  assign be_2x_13_30 = ~(px_13_30 & be_s2_13);
  assign be_2x_13_31 = ~(px_13_31 & be_s2_13);
  assign be_2x_13_32 = ~(px_13_32 & be_s2_13);
  assign be_2x_13_33 = ~(px_13_33 & be_s2_13);
  assign be_2x_13_4 = ~(px_13_4 & be_s2_13);
  assign be_2x_13_5 = ~(px_13_5 & be_s2_13);
  assign be_2x_13_6 = ~(px_13_6 & be_s2_13);
  assign be_2x_13_7 = ~(px_13_7 & be_s2_13);
  assign be_2x_13_8 = ~(px_13_8 & be_s2_13);
  assign be_2x_13_9 = ~(px_13_9 & be_s2_13);
  assign be_2x_14_0 = ~(px_14_0 & be_s2_14);
  assign be_2x_14_1 = ~(px_14_1 & be_s2_14);
  assign be_2x_14_10 = ~(px_14_10 & be_s2_14);
  assign be_2x_14_11 = ~(px_14_11 & be_s2_14);
  assign be_2x_14_12 = ~(px_14_12 & be_s2_14);
  assign be_2x_14_13 = ~(px_14_13 & be_s2_14);
  assign be_2x_14_14 = ~(px_14_14 & be_s2_14);
  assign be_2x_14_15 = ~(px_14_15 & be_s2_14);
  assign be_2x_14_16 = ~(px_14_16 & be_s2_14);
  assign be_2x_14_17 = ~(px_14_17 & be_s2_14);
  assign be_2x_14_18 = ~(px_14_18 & be_s2_14);
  assign be_2x_14_19 = ~(px_14_19 & be_s2_14);
  assign be_2x_14_2 = ~(px_14_2 & be_s2_14);
  assign be_2x_14_20 = ~(px_14_20 & be_s2_14);
  assign be_2x_14_21 = ~(px_14_21 & be_s2_14);
  assign be_2x_14_22 = ~(px_14_22 & be_s2_14);
  assign be_2x_14_23 = ~(px_14_23 & be_s2_14);
  assign be_2x_14_24 = ~(px_14_24 & be_s2_14);
  assign be_2x_14_25 = ~(px_14_25 & be_s2_14);
  assign be_2x_14_26 = ~(px_14_26 & be_s2_14);
  assign be_2x_14_27 = ~(px_14_27 & be_s2_14);
  assign be_2x_14_28 = ~(px_14_28 & be_s2_14);
  assign be_2x_14_29 = ~(px_14_29 & be_s2_14);
  assign be_2x_14_3 = ~(px_14_3 & be_s2_14);
  assign be_2x_14_30 = ~(px_14_30 & be_s2_14);
  assign be_2x_14_31 = ~(px_14_31 & be_s2_14);
  assign be_2x_14_32 = ~(px_14_32 & be_s2_14);
  assign be_2x_14_33 = ~(px_14_33 & be_s2_14);
  assign be_2x_14_4 = ~(px_14_4 & be_s2_14);
  assign be_2x_14_5 = ~(px_14_5 & be_s2_14);
  assign be_2x_14_6 = ~(px_14_6 & be_s2_14);
  assign be_2x_14_7 = ~(px_14_7 & be_s2_14);
  assign be_2x_14_8 = ~(px_14_8 & be_s2_14);
  assign be_2x_14_9 = ~(px_14_9 & be_s2_14);
  assign be_2x_15_0 = ~(px_15_0 & be_s2_15);
  assign be_2x_15_1 = ~(px_15_1 & be_s2_15);
  assign be_2x_15_10 = ~(px_15_10 & be_s2_15);
  assign be_2x_15_11 = ~(px_15_11 & be_s2_15);
  assign be_2x_15_12 = ~(px_15_12 & be_s2_15);
  assign be_2x_15_13 = ~(px_15_13 & be_s2_15);
  assign be_2x_15_14 = ~(px_15_14 & be_s2_15);
  assign be_2x_15_15 = ~(px_15_15 & be_s2_15);
  assign be_2x_15_16 = ~(px_15_16 & be_s2_15);
  assign be_2x_15_17 = ~(px_15_17 & be_s2_15);
  assign be_2x_15_18 = ~(px_15_18 & be_s2_15);
  assign be_2x_15_19 = ~(px_15_19 & be_s2_15);
  assign be_2x_15_2 = ~(px_15_2 & be_s2_15);
  assign be_2x_15_20 = ~(px_15_20 & be_s2_15);
  assign be_2x_15_21 = ~(px_15_21 & be_s2_15);
  assign be_2x_15_22 = ~(px_15_22 & be_s2_15);
  assign be_2x_15_23 = ~(px_15_23 & be_s2_15);
  assign be_2x_15_24 = ~(px_15_24 & be_s2_15);
  assign be_2x_15_25 = ~(px_15_25 & be_s2_15);
  assign be_2x_15_26 = ~(px_15_26 & be_s2_15);
  assign be_2x_15_27 = ~(px_15_27 & be_s2_15);
  assign be_2x_15_28 = ~(px_15_28 & be_s2_15);
  assign be_2x_15_29 = ~(px_15_29 & be_s2_15);
  assign be_2x_15_3 = ~(px_15_3 & be_s2_15);
  assign be_2x_15_30 = ~(px_15_30 & be_s2_15);
  assign be_2x_15_31 = ~(px_15_31 & be_s2_15);
  assign be_2x_15_32 = ~(px_15_32 & be_s2_15);
  assign be_2x_15_33 = ~(px_15_33 & be_s2_15);
  assign be_2x_15_4 = ~(px_15_4 & be_s2_15);
  assign be_2x_15_5 = ~(px_15_5 & be_s2_15);
  assign be_2x_15_6 = ~(px_15_6 & be_s2_15);
  assign be_2x_15_7 = ~(px_15_7 & be_s2_15);
  assign be_2x_15_8 = ~(px_15_8 & be_s2_15);
  assign be_2x_15_9 = ~(px_15_9 & be_s2_15);
  assign be_2x_16_0 = ~(px_16_0 & be_s2_16);
  assign be_2x_16_1 = ~(px_16_1 & be_s2_16);
  assign be_2x_16_10 = ~(px_16_10 & be_s2_16);
  assign be_2x_16_11 = ~(px_16_11 & be_s2_16);
  assign be_2x_16_12 = ~(px_16_12 & be_s2_16);
  assign be_2x_16_13 = ~(px_16_13 & be_s2_16);
  assign be_2x_16_14 = ~(px_16_14 & be_s2_16);
  assign be_2x_16_15 = ~(px_16_15 & be_s2_16);
  assign be_2x_16_16 = ~(px_16_16 & be_s2_16);
  assign be_2x_16_17 = ~(px_16_17 & be_s2_16);
  assign be_2x_16_18 = ~(px_16_18 & be_s2_16);
  assign be_2x_16_19 = ~(px_16_19 & be_s2_16);
  assign be_2x_16_2 = ~(px_16_2 & be_s2_16);
  assign be_2x_16_20 = ~(px_16_20 & be_s2_16);
  assign be_2x_16_21 = ~(px_16_21 & be_s2_16);
  assign be_2x_16_22 = ~(px_16_22 & be_s2_16);
  assign be_2x_16_23 = ~(px_16_23 & be_s2_16);
  assign be_2x_16_24 = ~(px_16_24 & be_s2_16);
  assign be_2x_16_25 = ~(px_16_25 & be_s2_16);
  assign be_2x_16_26 = ~(px_16_26 & be_s2_16);
  assign be_2x_16_27 = ~(px_16_27 & be_s2_16);
  assign be_2x_16_28 = ~(px_16_28 & be_s2_16);
  assign be_2x_16_29 = ~(px_16_29 & be_s2_16);
  assign be_2x_16_3 = ~(px_16_3 & be_s2_16);
  assign be_2x_16_30 = ~(px_16_30 & be_s2_16);
  assign be_2x_16_31 = ~(px_16_31 & be_s2_16);
  assign be_2x_16_4 = ~(px_16_4 & be_s2_16);
  assign be_2x_16_5 = ~(px_16_5 & be_s2_16);
  assign be_2x_16_6 = ~(px_16_6 & be_s2_16);
  assign be_2x_16_7 = ~(px_16_7 & be_s2_16);
  assign be_2x_16_8 = ~(px_16_8 & be_s2_16);
  assign be_2x_16_9 = ~(px_16_9 & be_s2_16);
  assign be_2x_1_0 = ~(px_1_0 & be_s2_1);
  assign be_2x_1_1 = ~(px_1_1 & be_s2_1);
  assign be_2x_1_10 = ~(px_1_10 & be_s2_1);
  assign be_2x_1_11 = ~(px_1_11 & be_s2_1);
  assign be_2x_1_12 = ~(px_1_12 & be_s2_1);
  assign be_2x_1_13 = ~(px_1_13 & be_s2_1);
  assign be_2x_1_14 = ~(px_1_14 & be_s2_1);
  assign be_2x_1_15 = ~(px_1_15 & be_s2_1);
  assign be_2x_1_16 = ~(px_1_16 & be_s2_1);
  assign be_2x_1_17 = ~(px_1_17 & be_s2_1);
  assign be_2x_1_18 = ~(px_1_18 & be_s2_1);
  assign be_2x_1_19 = ~(px_1_19 & be_s2_1);
  assign be_2x_1_2 = ~(px_1_2 & be_s2_1);
  assign be_2x_1_20 = ~(px_1_20 & be_s2_1);
  assign be_2x_1_21 = ~(px_1_21 & be_s2_1);
  assign be_2x_1_22 = ~(px_1_22 & be_s2_1);
  assign be_2x_1_23 = ~(px_1_23 & be_s2_1);
  assign be_2x_1_24 = ~(px_1_24 & be_s2_1);
  assign be_2x_1_25 = ~(px_1_25 & be_s2_1);
  assign be_2x_1_26 = ~(px_1_26 & be_s2_1);
  assign be_2x_1_27 = ~(px_1_27 & be_s2_1);
  assign be_2x_1_28 = ~(px_1_28 & be_s2_1);
  assign be_2x_1_29 = ~(px_1_29 & be_s2_1);
  assign be_2x_1_3 = ~(px_1_3 & be_s2_1);
  assign be_2x_1_30 = ~(px_1_30 & be_s2_1);
  assign be_2x_1_31 = ~(px_1_31 & be_s2_1);
  assign be_2x_1_32 = ~(px_1_32 & be_s2_1);
  assign be_2x_1_33 = ~(px_1_33 & be_s2_1);
  assign be_2x_1_4 = ~(px_1_4 & be_s2_1);
  assign be_2x_1_5 = ~(px_1_5 & be_s2_1);
  assign be_2x_1_6 = ~(px_1_6 & be_s2_1);
  assign be_2x_1_7 = ~(px_1_7 & be_s2_1);
  assign be_2x_1_8 = ~(px_1_8 & be_s2_1);
  assign be_2x_1_9 = ~(px_1_9 & be_s2_1);
  assign be_2x_2_0 = ~(px_2_0 & be_s2_2);
  assign be_2x_2_1 = ~(px_2_1 & be_s2_2);
  assign be_2x_2_10 = ~(px_2_10 & be_s2_2);
  assign be_2x_2_11 = ~(px_2_11 & be_s2_2);
  assign be_2x_2_12 = ~(px_2_12 & be_s2_2);
  assign be_2x_2_13 = ~(px_2_13 & be_s2_2);
  assign be_2x_2_14 = ~(px_2_14 & be_s2_2);
  assign be_2x_2_15 = ~(px_2_15 & be_s2_2);
  assign be_2x_2_16 = ~(px_2_16 & be_s2_2);
  assign be_2x_2_17 = ~(px_2_17 & be_s2_2);
  assign be_2x_2_18 = ~(px_2_18 & be_s2_2);
  assign be_2x_2_19 = ~(px_2_19 & be_s2_2);
  assign be_2x_2_2 = ~(px_2_2 & be_s2_2);
  assign be_2x_2_20 = ~(px_2_20 & be_s2_2);
  assign be_2x_2_21 = ~(px_2_21 & be_s2_2);
  assign be_2x_2_22 = ~(px_2_22 & be_s2_2);
  assign be_2x_2_23 = ~(px_2_23 & be_s2_2);
  assign be_2x_2_24 = ~(px_2_24 & be_s2_2);
  assign be_2x_2_25 = ~(px_2_25 & be_s2_2);
  assign be_2x_2_26 = ~(px_2_26 & be_s2_2);
  assign be_2x_2_27 = ~(px_2_27 & be_s2_2);
  assign be_2x_2_28 = ~(px_2_28 & be_s2_2);
  assign be_2x_2_29 = ~(px_2_29 & be_s2_2);
  assign be_2x_2_3 = ~(px_2_3 & be_s2_2);
  assign be_2x_2_30 = ~(px_2_30 & be_s2_2);
  assign be_2x_2_31 = ~(px_2_31 & be_s2_2);
  assign be_2x_2_32 = ~(px_2_32 & be_s2_2);
  assign be_2x_2_33 = ~(px_2_33 & be_s2_2);
  assign be_2x_2_4 = ~(px_2_4 & be_s2_2);
  assign be_2x_2_5 = ~(px_2_5 & be_s2_2);
  assign be_2x_2_6 = ~(px_2_6 & be_s2_2);
  assign be_2x_2_7 = ~(px_2_7 & be_s2_2);
  assign be_2x_2_8 = ~(px_2_8 & be_s2_2);
  assign be_2x_2_9 = ~(px_2_9 & be_s2_2);
  assign be_2x_3_0 = ~(px_3_0 & be_s2_3);
  assign be_2x_3_1 = ~(px_3_1 & be_s2_3);
  assign be_2x_3_10 = ~(px_3_10 & be_s2_3);
  assign be_2x_3_11 = ~(px_3_11 & be_s2_3);
  assign be_2x_3_12 = ~(px_3_12 & be_s2_3);
  assign be_2x_3_13 = ~(px_3_13 & be_s2_3);
  assign be_2x_3_14 = ~(px_3_14 & be_s2_3);
  assign be_2x_3_15 = ~(px_3_15 & be_s2_3);
  assign be_2x_3_16 = ~(px_3_16 & be_s2_3);
  assign be_2x_3_17 = ~(px_3_17 & be_s2_3);
  assign be_2x_3_18 = ~(px_3_18 & be_s2_3);
  assign be_2x_3_19 = ~(px_3_19 & be_s2_3);
  assign be_2x_3_2 = ~(px_3_2 & be_s2_3);
  assign be_2x_3_20 = ~(px_3_20 & be_s2_3);
  assign be_2x_3_21 = ~(px_3_21 & be_s2_3);
  assign be_2x_3_22 = ~(px_3_22 & be_s2_3);
  assign be_2x_3_23 = ~(px_3_23 & be_s2_3);
  assign be_2x_3_24 = ~(px_3_24 & be_s2_3);
  assign be_2x_3_25 = ~(px_3_25 & be_s2_3);
  assign be_2x_3_26 = ~(px_3_26 & be_s2_3);
  assign be_2x_3_27 = ~(px_3_27 & be_s2_3);
  assign be_2x_3_28 = ~(px_3_28 & be_s2_3);
  assign be_2x_3_29 = ~(px_3_29 & be_s2_3);
  assign be_2x_3_3 = ~(px_3_3 & be_s2_3);
  assign be_2x_3_30 = ~(px_3_30 & be_s2_3);
  assign be_2x_3_31 = ~(px_3_31 & be_s2_3);
  assign be_2x_3_32 = ~(px_3_32 & be_s2_3);
  assign be_2x_3_33 = ~(px_3_33 & be_s2_3);
  assign be_2x_3_4 = ~(px_3_4 & be_s2_3);
  assign be_2x_3_5 = ~(px_3_5 & be_s2_3);
  assign be_2x_3_6 = ~(px_3_6 & be_s2_3);
  assign be_2x_3_7 = ~(px_3_7 & be_s2_3);
  assign be_2x_3_8 = ~(px_3_8 & be_s2_3);
  assign be_2x_3_9 = ~(px_3_9 & be_s2_3);
  assign be_2x_4_0 = ~(px_4_0 & be_s2_4);
  assign be_2x_4_1 = ~(px_4_1 & be_s2_4);
  assign be_2x_4_10 = ~(px_4_10 & be_s2_4);
  assign be_2x_4_11 = ~(px_4_11 & be_s2_4);
  assign be_2x_4_12 = ~(px_4_12 & be_s2_4);
  assign be_2x_4_13 = ~(px_4_13 & be_s2_4);
  assign be_2x_4_14 = ~(px_4_14 & be_s2_4);
  assign be_2x_4_15 = ~(px_4_15 & be_s2_4);
  assign be_2x_4_16 = ~(px_4_16 & be_s2_4);
  assign be_2x_4_17 = ~(px_4_17 & be_s2_4);
  assign be_2x_4_18 = ~(px_4_18 & be_s2_4);
  assign be_2x_4_19 = ~(px_4_19 & be_s2_4);
  assign be_2x_4_2 = ~(px_4_2 & be_s2_4);
  assign be_2x_4_20 = ~(px_4_20 & be_s2_4);
  assign be_2x_4_21 = ~(px_4_21 & be_s2_4);
  assign be_2x_4_22 = ~(px_4_22 & be_s2_4);
  assign be_2x_4_23 = ~(px_4_23 & be_s2_4);
  assign be_2x_4_24 = ~(px_4_24 & be_s2_4);
  assign be_2x_4_25 = ~(px_4_25 & be_s2_4);
  assign be_2x_4_26 = ~(px_4_26 & be_s2_4);
  assign be_2x_4_27 = ~(px_4_27 & be_s2_4);
  assign be_2x_4_28 = ~(px_4_28 & be_s2_4);
  assign be_2x_4_29 = ~(px_4_29 & be_s2_4);
  assign be_2x_4_3 = ~(px_4_3 & be_s2_4);
  assign be_2x_4_30 = ~(px_4_30 & be_s2_4);
  assign be_2x_4_31 = ~(px_4_31 & be_s2_4);
  assign be_2x_4_32 = ~(px_4_32 & be_s2_4);
  assign be_2x_4_33 = ~(px_4_33 & be_s2_4);
  assign be_2x_4_4 = ~(px_4_4 & be_s2_4);
  assign be_2x_4_5 = ~(px_4_5 & be_s2_4);
  assign be_2x_4_6 = ~(px_4_6 & be_s2_4);
  assign be_2x_4_7 = ~(px_4_7 & be_s2_4);
  assign be_2x_4_8 = ~(px_4_8 & be_s2_4);
  assign be_2x_4_9 = ~(px_4_9 & be_s2_4);
  assign be_2x_5_0 = ~(px_5_0 & be_s2_5);
  assign be_2x_5_1 = ~(px_5_1 & be_s2_5);
  assign be_2x_5_10 = ~(px_5_10 & be_s2_5);
  assign be_2x_5_11 = ~(px_5_11 & be_s2_5);
  assign be_2x_5_12 = ~(px_5_12 & be_s2_5);
  assign be_2x_5_13 = ~(px_5_13 & be_s2_5);
  assign be_2x_5_14 = ~(px_5_14 & be_s2_5);
  assign be_2x_5_15 = ~(px_5_15 & be_s2_5);
  assign be_2x_5_16 = ~(px_5_16 & be_s2_5);
  assign be_2x_5_17 = ~(px_5_17 & be_s2_5);
  assign be_2x_5_18 = ~(px_5_18 & be_s2_5);
  assign be_2x_5_19 = ~(px_5_19 & be_s2_5);
  assign be_2x_5_2 = ~(px_5_2 & be_s2_5);
  assign be_2x_5_20 = ~(px_5_20 & be_s2_5);
  assign be_2x_5_21 = ~(px_5_21 & be_s2_5);
  assign be_2x_5_22 = ~(px_5_22 & be_s2_5);
  assign be_2x_5_23 = ~(px_5_23 & be_s2_5);
  assign be_2x_5_24 = ~(px_5_24 & be_s2_5);
  assign be_2x_5_25 = ~(px_5_25 & be_s2_5);
  assign be_2x_5_26 = ~(px_5_26 & be_s2_5);
  assign be_2x_5_27 = ~(px_5_27 & be_s2_5);
  assign be_2x_5_28 = ~(px_5_28 & be_s2_5);
  assign be_2x_5_29 = ~(px_5_29 & be_s2_5);
  assign be_2x_5_3 = ~(px_5_3 & be_s2_5);
  assign be_2x_5_30 = ~(px_5_30 & be_s2_5);
  assign be_2x_5_31 = ~(px_5_31 & be_s2_5);
  assign be_2x_5_32 = ~(px_5_32 & be_s2_5);
  assign be_2x_5_33 = ~(px_5_33 & be_s2_5);
  assign be_2x_5_4 = ~(px_5_4 & be_s2_5);
  assign be_2x_5_5 = ~(px_5_5 & be_s2_5);
  assign be_2x_5_6 = ~(px_5_6 & be_s2_5);
  assign be_2x_5_7 = ~(px_5_7 & be_s2_5);
  assign be_2x_5_8 = ~(px_5_8 & be_s2_5);
  assign be_2x_5_9 = ~(px_5_9 & be_s2_5);
  assign be_2x_6_0 = ~(px_6_0 & be_s2_6);
  assign be_2x_6_1 = ~(px_6_1 & be_s2_6);
  assign be_2x_6_10 = ~(px_6_10 & be_s2_6);
  assign be_2x_6_11 = ~(px_6_11 & be_s2_6);
  assign be_2x_6_12 = ~(px_6_12 & be_s2_6);
  assign be_2x_6_13 = ~(px_6_13 & be_s2_6);
  assign be_2x_6_14 = ~(px_6_14 & be_s2_6);
  assign be_2x_6_15 = ~(px_6_15 & be_s2_6);
  assign be_2x_6_16 = ~(px_6_16 & be_s2_6);
  assign be_2x_6_17 = ~(px_6_17 & be_s2_6);
  assign be_2x_6_18 = ~(px_6_18 & be_s2_6);
  assign be_2x_6_19 = ~(px_6_19 & be_s2_6);
  assign be_2x_6_2 = ~(px_6_2 & be_s2_6);
  assign be_2x_6_20 = ~(px_6_20 & be_s2_6);
  assign be_2x_6_21 = ~(px_6_21 & be_s2_6);
  assign be_2x_6_22 = ~(px_6_22 & be_s2_6);
  assign be_2x_6_23 = ~(px_6_23 & be_s2_6);
  assign be_2x_6_24 = ~(px_6_24 & be_s2_6);
  assign be_2x_6_25 = ~(px_6_25 & be_s2_6);
  assign be_2x_6_26 = ~(px_6_26 & be_s2_6);
  assign be_2x_6_27 = ~(px_6_27 & be_s2_6);
  assign be_2x_6_28 = ~(px_6_28 & be_s2_6);
  assign be_2x_6_29 = ~(px_6_29 & be_s2_6);
  assign be_2x_6_3 = ~(px_6_3 & be_s2_6);
  assign be_2x_6_30 = ~(px_6_30 & be_s2_6);
  assign be_2x_6_31 = ~(px_6_31 & be_s2_6);
  assign be_2x_6_32 = ~(px_6_32 & be_s2_6);
  assign be_2x_6_33 = ~(px_6_33 & be_s2_6);
  assign be_2x_6_4 = ~(px_6_4 & be_s2_6);
  assign be_2x_6_5 = ~(px_6_5 & be_s2_6);
  assign be_2x_6_6 = ~(px_6_6 & be_s2_6);
  assign be_2x_6_7 = ~(px_6_7 & be_s2_6);
  assign be_2x_6_8 = ~(px_6_8 & be_s2_6);
  assign be_2x_6_9 = ~(px_6_9 & be_s2_6);
  assign be_2x_7_0 = ~(px_7_0 & be_s2_7);
  assign be_2x_7_1 = ~(px_7_1 & be_s2_7);
  assign be_2x_7_10 = ~(px_7_10 & be_s2_7);
  assign be_2x_7_11 = ~(px_7_11 & be_s2_7);
  assign be_2x_7_12 = ~(px_7_12 & be_s2_7);
  assign be_2x_7_13 = ~(px_7_13 & be_s2_7);
  assign be_2x_7_14 = ~(px_7_14 & be_s2_7);
  assign be_2x_7_15 = ~(px_7_15 & be_s2_7);
  assign be_2x_7_16 = ~(px_7_16 & be_s2_7);
  assign be_2x_7_17 = ~(px_7_17 & be_s2_7);
  assign be_2x_7_18 = ~(px_7_18 & be_s2_7);
  assign be_2x_7_19 = ~(px_7_19 & be_s2_7);
  assign be_2x_7_2 = ~(px_7_2 & be_s2_7);
  assign be_2x_7_20 = ~(px_7_20 & be_s2_7);
  assign be_2x_7_21 = ~(px_7_21 & be_s2_7);
  assign be_2x_7_22 = ~(px_7_22 & be_s2_7);
  assign be_2x_7_23 = ~(px_7_23 & be_s2_7);
  assign be_2x_7_24 = ~(px_7_24 & be_s2_7);
  assign be_2x_7_25 = ~(px_7_25 & be_s2_7);
  assign be_2x_7_26 = ~(px_7_26 & be_s2_7);
  assign be_2x_7_27 = ~(px_7_27 & be_s2_7);
  assign be_2x_7_28 = ~(px_7_28 & be_s2_7);
  assign be_2x_7_29 = ~(px_7_29 & be_s2_7);
  assign be_2x_7_3 = ~(px_7_3 & be_s2_7);
  assign be_2x_7_30 = ~(px_7_30 & be_s2_7);
  assign be_2x_7_31 = ~(px_7_31 & be_s2_7);
  assign be_2x_7_32 = ~(px_7_32 & be_s2_7);
  assign be_2x_7_33 = ~(px_7_33 & be_s2_7);
  assign be_2x_7_4 = ~(px_7_4 & be_s2_7);
  assign be_2x_7_5 = ~(px_7_5 & be_s2_7);
  assign be_2x_7_6 = ~(px_7_6 & be_s2_7);
  assign be_2x_7_7 = ~(px_7_7 & be_s2_7);
  assign be_2x_7_8 = ~(px_7_8 & be_s2_7);
  assign be_2x_7_9 = ~(px_7_9 & be_s2_7);
  assign be_2x_8_0 = ~(px_8_0 & be_s2_8);
  assign be_2x_8_1 = ~(px_8_1 & be_s2_8);
  assign be_2x_8_10 = ~(px_8_10 & be_s2_8);
  assign be_2x_8_11 = ~(px_8_11 & be_s2_8);
  assign be_2x_8_12 = ~(px_8_12 & be_s2_8);
  assign be_2x_8_13 = ~(px_8_13 & be_s2_8);
  assign be_2x_8_14 = ~(px_8_14 & be_s2_8);
  assign be_2x_8_15 = ~(px_8_15 & be_s2_8);
  assign be_2x_8_16 = ~(px_8_16 & be_s2_8);
  assign be_2x_8_17 = ~(px_8_17 & be_s2_8);
  assign be_2x_8_18 = ~(px_8_18 & be_s2_8);
  assign be_2x_8_19 = ~(px_8_19 & be_s2_8);
  assign be_2x_8_2 = ~(px_8_2 & be_s2_8);
  assign be_2x_8_20 = ~(px_8_20 & be_s2_8);
  assign be_2x_8_21 = ~(px_8_21 & be_s2_8);
  assign be_2x_8_22 = ~(px_8_22 & be_s2_8);
  assign be_2x_8_23 = ~(px_8_23 & be_s2_8);
  assign be_2x_8_24 = ~(px_8_24 & be_s2_8);
  assign be_2x_8_25 = ~(px_8_25 & be_s2_8);
  assign be_2x_8_26 = ~(px_8_26 & be_s2_8);
  assign be_2x_8_27 = ~(px_8_27 & be_s2_8);
  assign be_2x_8_28 = ~(px_8_28 & be_s2_8);
  assign be_2x_8_29 = ~(px_8_29 & be_s2_8);
  assign be_2x_8_3 = ~(px_8_3 & be_s2_8);
  assign be_2x_8_30 = ~(px_8_30 & be_s2_8);
  assign be_2x_8_31 = ~(px_8_31 & be_s2_8);
  assign be_2x_8_32 = ~(px_8_32 & be_s2_8);
  assign be_2x_8_33 = ~(px_8_33 & be_s2_8);
  assign be_2x_8_4 = ~(px_8_4 & be_s2_8);
  assign be_2x_8_5 = ~(px_8_5 & be_s2_8);
  assign be_2x_8_6 = ~(px_8_6 & be_s2_8);
  assign be_2x_8_7 = ~(px_8_7 & be_s2_8);
  assign be_2x_8_8 = ~(px_8_8 & be_s2_8);
  assign be_2x_8_9 = ~(px_8_9 & be_s2_8);
  assign be_2x_9_0 = ~(px_9_0 & be_s2_9);
  assign be_2x_9_1 = ~(px_9_1 & be_s2_9);
  assign be_2x_9_10 = ~(px_9_10 & be_s2_9);
  assign be_2x_9_11 = ~(px_9_11 & be_s2_9);
  assign be_2x_9_12 = ~(px_9_12 & be_s2_9);
  assign be_2x_9_13 = ~(px_9_13 & be_s2_9);
  assign be_2x_9_14 = ~(px_9_14 & be_s2_9);
  assign be_2x_9_15 = ~(px_9_15 & be_s2_9);
  assign be_2x_9_16 = ~(px_9_16 & be_s2_9);
  assign be_2x_9_17 = ~(px_9_17 & be_s2_9);
  assign be_2x_9_18 = ~(px_9_18 & be_s2_9);
  assign be_2x_9_19 = ~(px_9_19 & be_s2_9);
  assign be_2x_9_2 = ~(px_9_2 & be_s2_9);
  assign be_2x_9_20 = ~(px_9_20 & be_s2_9);
  assign be_2x_9_21 = ~(px_9_21 & be_s2_9);
  assign be_2x_9_22 = ~(px_9_22 & be_s2_9);
  assign be_2x_9_23 = ~(px_9_23 & be_s2_9);
  assign be_2x_9_24 = ~(px_9_24 & be_s2_9);
  assign be_2x_9_25 = ~(px_9_25 & be_s2_9);
  assign be_2x_9_26 = ~(px_9_26 & be_s2_9);
  assign be_2x_9_27 = ~(px_9_27 & be_s2_9);
  assign be_2x_9_28 = ~(px_9_28 & be_s2_9);
  assign be_2x_9_29 = ~(px_9_29 & be_s2_9);
  assign be_2x_9_3 = ~(px_9_3 & be_s2_9);
  assign be_2x_9_30 = ~(px_9_30 & be_s2_9);
  assign be_2x_9_31 = ~(px_9_31 & be_s2_9);
  assign be_2x_9_32 = ~(px_9_32 & be_s2_9);
  assign be_2x_9_33 = ~(px_9_33 & be_s2_9);
  assign be_2x_9_4 = ~(px_9_4 & be_s2_9);
  assign be_2x_9_5 = ~(px_9_5 & be_s2_9);
  assign be_2x_9_6 = ~(px_9_6 & be_s2_9);
  assign be_2x_9_7 = ~(px_9_7 & be_s2_9);
  assign be_2x_9_8 = ~(px_9_8 & be_s2_9);
  assign be_2x_9_9 = ~(px_9_9 & be_s2_9);
  assign be_c_0 = be_d_0 & be_neg_0;
  assign be_c_1 = be_d_1 & be_neg_1;
  assign be_c_10 = be_d_10 & be_neg_10;
  assign be_c_11 = be_d_11 & be_neg_11;
  assign be_c_12 = be_d_12 & be_neg_12;
  assign be_c_13 = be_d_13 & be_neg_13;
  assign be_c_14 = be_d_14 & be_neg_14;
  assign be_c_15 = be_d_15 & be_neg_15;
  assign be_c_16 = be_d_16 & be_neg_16;
  assign be_c_2 = be_d_2 & be_neg_2;
  assign be_c_3 = be_d_3 & be_neg_3;
  assign be_c_4 = be_d_4 & be_neg_4;
  assign be_c_5 = be_d_5 & be_neg_5;
  assign be_c_6 = be_d_6 & be_neg_6;
  assign be_c_7 = be_d_7 & be_neg_7;
  assign be_c_8 = be_d_8 & be_neg_8;
  assign be_c_9 = be_d_9 & be_neg_9;
  assign be_d_0 = ny_0 | one;
  assign be_d_1 = ny_2 | ny_1;
  assign be_d_10 = ny_20 | ny_19;
  assign be_d_11 = ny_22 | ny_21;
  assign be_d_12 = ny_24 | ny_23;
  assign be_d_13 = ny_26 | ny_25;
  assign be_d_14 = ny_28 | ny_27;
  assign be_d_15 = ny_30 | ny_29;
  assign be_d_16 = one | ny_31;
  assign be_d_2 = ny_4 | ny_3;
  assign be_d_3 = ny_6 | ny_5;
  assign be_d_4 = ny_8 | ny_7;
  assign be_d_5 = ny_10 | ny_9;
  assign be_d_6 = ny_12 | ny_11;
  assign be_d_7 = ny_14 | ny_13;
  assign be_d_8 = ny_16 | ny_15;
  assign be_d_9 = ny_18 | ny_17;
  assign be_neg_0 = y_1;
  assign be_neg_1 = y_3;
  assign be_neg_10 = y_21;
  assign be_neg_11 = y_23;
  assign be_neg_12 = y_25;
  assign be_neg_13 = y_27;
  assign be_neg_14 = y_29;
  assign be_neg_15 = y_31;
  assign be_neg_16 = zero;
  assign be_neg_2 = y_5;
  assign be_neg_3 = y_7;
  assign be_neg_4 = y_9;
  assign be_neg_5 = y_11;
  assign be_neg_6 = y_13;
  assign be_neg_7 = y_15;
  assign be_neg_8 = y_17;
  assign be_neg_9 = y_19;
  assign be_s1_0 = y_0 ^ zero;
  assign be_s1_1 = y_2 ^ y_1;
  assign be_s1_10 = y_20 ^ y_19;
  assign be_s1_11 = y_22 ^ y_21;
  assign be_s1_12 = y_24 ^ y_23;
  assign be_s1_13 = y_26 ^ y_25;
  assign be_s1_14 = y_28 ^ y_27;
  assign be_s1_15 = y_30 ^ y_29;
  assign be_s1_16 = zero ^ y_31;
  assign be_s1_2 = y_4 ^ y_3;
  assign be_s1_3 = y_6 ^ y_5;
  assign be_s1_4 = y_8 ^ y_7;
  assign be_s1_5 = y_10 ^ y_9;
  assign be_s1_6 = y_12 ^ y_11;
  assign be_s1_7 = y_14 ^ y_13;
  assign be_s1_8 = y_16 ^ y_15;
  assign be_s1_9 = y_18 ^ y_17;
  assign be_s2_0 = be_s2_a_0 | be_s2_b_0;
  assign be_s2_1 = be_s2_a_1 | be_s2_b_1;
  assign be_s2_10 = be_s2_a_10 | be_s2_b_10;
  assign be_s2_11 = be_s2_a_11 | be_s2_b_11;
  assign be_s2_12 = be_s2_a_12 | be_s2_b_12;
  assign be_s2_13 = be_s2_a_13 | be_s2_b_13;
  assign be_s2_14 = be_s2_a_14 | be_s2_b_14;
  assign be_s2_15 = be_s2_a_15 | be_s2_b_15;
  assign be_s2_16 = be_s2_a_16 | be_s2_b_16;
  assign be_s2_2 = be_s2_a_2 | be_s2_b_2;
  assign be_s2_3 = be_s2_a_3 | be_s2_b_3;
  assign be_s2_4 = be_s2_a_4 | be_s2_b_4;
  assign be_s2_5 = be_s2_a_5 | be_s2_b_5;
  assign be_s2_6 = be_s2_a_6 | be_s2_b_6;
  assign be_s2_7 = be_s2_a_7 | be_s2_b_7;
  assign be_s2_8 = be_s2_a_8 | be_s2_b_8;
  assign be_s2_9 = be_s2_a_9 | be_s2_b_9;
  assign be_s2_a_0 = ny_1 & y_0 & zero;
  assign be_s2_a_1 = ny_3 & y_2 & y_1;
  assign be_s2_a_10 = ny_21 & y_20 & y_19;
  assign be_s2_a_11 = ny_23 & y_22 & y_21;
  assign be_s2_a_12 = ny_25 & y_24 & y_23;
  assign be_s2_a_13 = ny_27 & y_26 & y_25;
  assign be_s2_a_14 = ny_29 & y_28 & y_27;
  assign be_s2_a_15 = ny_31 & y_30 & y_29;
  assign be_s2_a_16 = one & zero & y_31;
  assign be_s2_a_2 = ny_5 & y_4 & y_3;
  assign be_s2_a_3 = ny_7 & y_6 & y_5;
  assign be_s2_a_4 = ny_9 & y_8 & y_7;
  assign be_s2_a_5 = ny_11 & y_10 & y_9;
  assign be_s2_a_6 = ny_13 & y_12 & y_11;
  assign be_s2_a_7 = ny_15 & y_14 & y_13;
  assign be_s2_a_8 = ny_17 & y_16 & y_15;
  assign be_s2_a_9 = ny_19 & y_18 & y_17;
  assign be_s2_b_0 = y_1 & ny_0 & one;
  assign be_s2_b_1 = y_3 & ny_2 & ny_1;
  assign be_s2_b_10 = y_21 & ny_20 & ny_19;
  assign be_s2_b_11 = y_23 & ny_22 & ny_21;
  assign be_s2_b_12 = y_25 & ny_24 & ny_23;
  assign be_s2_b_13 = y_27 & ny_26 & ny_25;
  assign be_s2_b_14 = y_29 & ny_28 & ny_27;
  assign be_s2_b_15 = y_31 & ny_30 & ny_29;
  assign be_s2_b_16 = zero & one & ny_31;
  assign be_s2_b_2 = y_5 & ny_4 & ny_3;
  assign be_s2_b_3 = y_7 & ny_6 & ny_5;
  assign be_s2_b_4 = y_9 & ny_8 & ny_7;
  assign be_s2_b_5 = y_11 & ny_10 & ny_9;
  assign be_s2_b_6 = y_13 & ny_12 & ny_11;
  assign be_s2_b_7 = y_15 & ny_14 & ny_13;
  assign be_s2_b_8 = y_17 & ny_16 & ny_15;
  assign be_s2_b_9 = y_19 & ny_18 & ny_17;
  assign be_x_0_0 = ~(px_0_1 & be_s1_0);
  assign be_x_0_1 = ~(px_0_2 & be_s1_0);
  assign be_x_0_10 = ~(px_0_11 & be_s1_0);
  assign be_x_0_11 = ~(px_0_12 & be_s1_0);
  assign be_x_0_12 = ~(px_0_13 & be_s1_0);
  assign be_x_0_13 = ~(px_0_14 & be_s1_0);
  assign be_x_0_14 = ~(px_0_15 & be_s1_0);
  assign be_x_0_15 = ~(px_0_16 & be_s1_0);
  assign be_x_0_16 = ~(px_0_17 & be_s1_0);
  assign be_x_0_17 = ~(px_0_18 & be_s1_0);
  assign be_x_0_18 = ~(px_0_19 & be_s1_0);
  assign be_x_0_19 = ~(px_0_20 & be_s1_0);
  assign be_x_0_2 = ~(px_0_3 & be_s1_0);
  assign be_x_0_20 = ~(px_0_21 & be_s1_0);
  assign be_x_0_21 = ~(px_0_22 & be_s1_0);
  assign be_x_0_22 = ~(px_0_23 & be_s1_0);
  assign be_x_0_23 = ~(px_0_24 & be_s1_0);
  assign be_x_0_24 = ~(px_0_25 & be_s1_0);
  assign be_x_0_25 = ~(px_0_26 & be_s1_0);
  assign be_x_0_26 = ~(px_0_27 & be_s1_0);
  assign be_x_0_27 = ~(px_0_28 & be_s1_0);
  assign be_x_0_28 = ~(px_0_29 & be_s1_0);
  assign be_x_0_29 = ~(px_0_30 & be_s1_0);
  assign be_x_0_3 = ~(px_0_4 & be_s1_0);
  assign be_x_0_30 = ~(px_0_31 & be_s1_0);
  assign be_x_0_31 = ~(px_0_32 & be_s1_0);
  assign be_x_0_32 = ~(px_0_33 & be_s1_0);
  assign be_x_0_33 = ~(px_0_34 & be_s1_0);
  assign be_x_0_4 = ~(px_0_5 & be_s1_0);
  assign be_x_0_5 = ~(px_0_6 & be_s1_0);
  assign be_x_0_6 = ~(px_0_7 & be_s1_0);
  assign be_x_0_7 = ~(px_0_8 & be_s1_0);
  assign be_x_0_8 = ~(px_0_9 & be_s1_0);
  assign be_x_0_9 = ~(px_0_10 & be_s1_0);
  assign be_x_10_0 = ~(px_10_1 & be_s1_10);
  assign be_x_10_1 = ~(px_10_2 & be_s1_10);
  assign be_x_10_10 = ~(px_10_11 & be_s1_10);
  assign be_x_10_11 = ~(px_10_12 & be_s1_10);
  assign be_x_10_12 = ~(px_10_13 & be_s1_10);
  assign be_x_10_13 = ~(px_10_14 & be_s1_10);
  assign be_x_10_14 = ~(px_10_15 & be_s1_10);
  assign be_x_10_15 = ~(px_10_16 & be_s1_10);
  assign be_x_10_16 = ~(px_10_17 & be_s1_10);
  assign be_x_10_17 = ~(px_10_18 & be_s1_10);
  assign be_x_10_18 = ~(px_10_19 & be_s1_10);
  assign be_x_10_19 = ~(px_10_20 & be_s1_10);
  assign be_x_10_2 = ~(px_10_3 & be_s1_10);
  assign be_x_10_20 = ~(px_10_21 & be_s1_10);
  assign be_x_10_21 = ~(px_10_22 & be_s1_10);
  assign be_x_10_22 = ~(px_10_23 & be_s1_10);
  assign be_x_10_23 = ~(px_10_24 & be_s1_10);
  assign be_x_10_24 = ~(px_10_25 & be_s1_10);
  assign be_x_10_25 = ~(px_10_26 & be_s1_10);
  assign be_x_10_26 = ~(px_10_27 & be_s1_10);
  assign be_x_10_27 = ~(px_10_28 & be_s1_10);
  assign be_x_10_28 = ~(px_10_29 & be_s1_10);
  assign be_x_10_29 = ~(px_10_30 & be_s1_10);
  assign be_x_10_3 = ~(px_10_4 & be_s1_10);
  assign be_x_10_30 = ~(px_10_31 & be_s1_10);
  assign be_x_10_31 = ~(px_10_32 & be_s1_10);
  assign be_x_10_32 = ~(px_10_33 & be_s1_10);
  assign be_x_10_33 = ~(px_10_34 & be_s1_10);
  assign be_x_10_4 = ~(px_10_5 & be_s1_10);
  assign be_x_10_5 = ~(px_10_6 & be_s1_10);
  assign be_x_10_6 = ~(px_10_7 & be_s1_10);
  assign be_x_10_7 = ~(px_10_8 & be_s1_10);
  assign be_x_10_8 = ~(px_10_9 & be_s1_10);
  assign be_x_10_9 = ~(px_10_10 & be_s1_10);
  assign be_x_11_0 = ~(px_11_1 & be_s1_11);
  assign be_x_11_1 = ~(px_11_2 & be_s1_11);
  assign be_x_11_10 = ~(px_11_11 & be_s1_11);
  assign be_x_11_11 = ~(px_11_12 & be_s1_11);
  assign be_x_11_12 = ~(px_11_13 & be_s1_11);
  assign be_x_11_13 = ~(px_11_14 & be_s1_11);
  assign be_x_11_14 = ~(px_11_15 & be_s1_11);
  assign be_x_11_15 = ~(px_11_16 & be_s1_11);
  assign be_x_11_16 = ~(px_11_17 & be_s1_11);
  assign be_x_11_17 = ~(px_11_18 & be_s1_11);
  assign be_x_11_18 = ~(px_11_19 & be_s1_11);
  assign be_x_11_19 = ~(px_11_20 & be_s1_11);
  assign be_x_11_2 = ~(px_11_3 & be_s1_11);
  assign be_x_11_20 = ~(px_11_21 & be_s1_11);
  assign be_x_11_21 = ~(px_11_22 & be_s1_11);
  assign be_x_11_22 = ~(px_11_23 & be_s1_11);
  assign be_x_11_23 = ~(px_11_24 & be_s1_11);
  assign be_x_11_24 = ~(px_11_25 & be_s1_11);
  assign be_x_11_25 = ~(px_11_26 & be_s1_11);
  assign be_x_11_26 = ~(px_11_27 & be_s1_11);
  assign be_x_11_27 = ~(px_11_28 & be_s1_11);
  assign be_x_11_28 = ~(px_11_29 & be_s1_11);
  assign be_x_11_29 = ~(px_11_30 & be_s1_11);
  assign be_x_11_3 = ~(px_11_4 & be_s1_11);
  assign be_x_11_30 = ~(px_11_31 & be_s1_11);
  assign be_x_11_31 = ~(px_11_32 & be_s1_11);
  assign be_x_11_32 = ~(px_11_33 & be_s1_11);
  assign be_x_11_33 = ~(px_11_34 & be_s1_11);
  assign be_x_11_4 = ~(px_11_5 & be_s1_11);
  assign be_x_11_5 = ~(px_11_6 & be_s1_11);
  assign be_x_11_6 = ~(px_11_7 & be_s1_11);
  assign be_x_11_7 = ~(px_11_8 & be_s1_11);
  assign be_x_11_8 = ~(px_11_9 & be_s1_11);
  assign be_x_11_9 = ~(px_11_10 & be_s1_11);
  assign be_x_12_0 = ~(px_12_1 & be_s1_12);
  assign be_x_12_1 = ~(px_12_2 & be_s1_12);
  assign be_x_12_10 = ~(px_12_11 & be_s1_12);
  assign be_x_12_11 = ~(px_12_12 & be_s1_12);
  assign be_x_12_12 = ~(px_12_13 & be_s1_12);
  assign be_x_12_13 = ~(px_12_14 & be_s1_12);
  assign be_x_12_14 = ~(px_12_15 & be_s1_12);
  assign be_x_12_15 = ~(px_12_16 & be_s1_12);
  assign be_x_12_16 = ~(px_12_17 & be_s1_12);
  assign be_x_12_17 = ~(px_12_18 & be_s1_12);
  assign be_x_12_18 = ~(px_12_19 & be_s1_12);
  assign be_x_12_19 = ~(px_12_20 & be_s1_12);
  assign be_x_12_2 = ~(px_12_3 & be_s1_12);
  assign be_x_12_20 = ~(px_12_21 & be_s1_12);
  assign be_x_12_21 = ~(px_12_22 & be_s1_12);
  assign be_x_12_22 = ~(px_12_23 & be_s1_12);
  assign be_x_12_23 = ~(px_12_24 & be_s1_12);
  assign be_x_12_24 = ~(px_12_25 & be_s1_12);
  assign be_x_12_25 = ~(px_12_26 & be_s1_12);
  assign be_x_12_26 = ~(px_12_27 & be_s1_12);
  assign be_x_12_27 = ~(px_12_28 & be_s1_12);
  assign be_x_12_28 = ~(px_12_29 & be_s1_12);
  assign be_x_12_29 = ~(px_12_30 & be_s1_12);
  assign be_x_12_3 = ~(px_12_4 & be_s1_12);
  assign be_x_12_30 = ~(px_12_31 & be_s1_12);
  assign be_x_12_31 = ~(px_12_32 & be_s1_12);
  assign be_x_12_32 = ~(px_12_33 & be_s1_12);
  assign be_x_12_33 = ~(px_12_34 & be_s1_12);
  assign be_x_12_4 = ~(px_12_5 & be_s1_12);
  assign be_x_12_5 = ~(px_12_6 & be_s1_12);
  assign be_x_12_6 = ~(px_12_7 & be_s1_12);
  assign be_x_12_7 = ~(px_12_8 & be_s1_12);
  assign be_x_12_8 = ~(px_12_9 & be_s1_12);
  assign be_x_12_9 = ~(px_12_10 & be_s1_12);
  assign be_x_13_0 = ~(px_13_1 & be_s1_13);
  assign be_x_13_1 = ~(px_13_2 & be_s1_13);
  assign be_x_13_10 = ~(px_13_11 & be_s1_13);
  assign be_x_13_11 = ~(px_13_12 & be_s1_13);
  assign be_x_13_12 = ~(px_13_13 & be_s1_13);
  assign be_x_13_13 = ~(px_13_14 & be_s1_13);
  assign be_x_13_14 = ~(px_13_15 & be_s1_13);
  assign be_x_13_15 = ~(px_13_16 & be_s1_13);
  assign be_x_13_16 = ~(px_13_17 & be_s1_13);
  assign be_x_13_17 = ~(px_13_18 & be_s1_13);
  assign be_x_13_18 = ~(px_13_19 & be_s1_13);
  assign be_x_13_19 = ~(px_13_20 & be_s1_13);
  assign be_x_13_2 = ~(px_13_3 & be_s1_13);
  assign be_x_13_20 = ~(px_13_21 & be_s1_13);
  assign be_x_13_21 = ~(px_13_22 & be_s1_13);
  assign be_x_13_22 = ~(px_13_23 & be_s1_13);
  assign be_x_13_23 = ~(px_13_24 & be_s1_13);
  assign be_x_13_24 = ~(px_13_25 & be_s1_13);
  assign be_x_13_25 = ~(px_13_26 & be_s1_13);
  assign be_x_13_26 = ~(px_13_27 & be_s1_13);
  assign be_x_13_27 = ~(px_13_28 & be_s1_13);
  assign be_x_13_28 = ~(px_13_29 & be_s1_13);
  assign be_x_13_29 = ~(px_13_30 & be_s1_13);
  assign be_x_13_3 = ~(px_13_4 & be_s1_13);
  assign be_x_13_30 = ~(px_13_31 & be_s1_13);
  assign be_x_13_31 = ~(px_13_32 & be_s1_13);
  assign be_x_13_32 = ~(px_13_33 & be_s1_13);
  assign be_x_13_33 = ~(px_13_34 & be_s1_13);
  assign be_x_13_4 = ~(px_13_5 & be_s1_13);
  assign be_x_13_5 = ~(px_13_6 & be_s1_13);
  assign be_x_13_6 = ~(px_13_7 & be_s1_13);
  assign be_x_13_7 = ~(px_13_8 & be_s1_13);
  assign be_x_13_8 = ~(px_13_9 & be_s1_13);
  assign be_x_13_9 = ~(px_13_10 & be_s1_13);
  assign be_x_14_0 = ~(px_14_1 & be_s1_14);
  assign be_x_14_1 = ~(px_14_2 & be_s1_14);
  assign be_x_14_10 = ~(px_14_11 & be_s1_14);
  assign be_x_14_11 = ~(px_14_12 & be_s1_14);
  assign be_x_14_12 = ~(px_14_13 & be_s1_14);
  assign be_x_14_13 = ~(px_14_14 & be_s1_14);
  assign be_x_14_14 = ~(px_14_15 & be_s1_14);
  assign be_x_14_15 = ~(px_14_16 & be_s1_14);
  assign be_x_14_16 = ~(px_14_17 & be_s1_14);
  assign be_x_14_17 = ~(px_14_18 & be_s1_14);
  assign be_x_14_18 = ~(px_14_19 & be_s1_14);
  assign be_x_14_19 = ~(px_14_20 & be_s1_14);
  assign be_x_14_2 = ~(px_14_3 & be_s1_14);
  assign be_x_14_20 = ~(px_14_21 & be_s1_14);
  assign be_x_14_21 = ~(px_14_22 & be_s1_14);
  assign be_x_14_22 = ~(px_14_23 & be_s1_14);
  assign be_x_14_23 = ~(px_14_24 & be_s1_14);
  assign be_x_14_24 = ~(px_14_25 & be_s1_14);
  assign be_x_14_25 = ~(px_14_26 & be_s1_14);
  assign be_x_14_26 = ~(px_14_27 & be_s1_14);
  assign be_x_14_27 = ~(px_14_28 & be_s1_14);
  assign be_x_14_28 = ~(px_14_29 & be_s1_14);
  assign be_x_14_29 = ~(px_14_30 & be_s1_14);
  assign be_x_14_3 = ~(px_14_4 & be_s1_14);
  assign be_x_14_30 = ~(px_14_31 & be_s1_14);
  assign be_x_14_31 = ~(px_14_32 & be_s1_14);
  assign be_x_14_32 = ~(px_14_33 & be_s1_14);
  assign be_x_14_33 = ~(px_14_34 & be_s1_14);
  assign be_x_14_4 = ~(px_14_5 & be_s1_14);
  assign be_x_14_5 = ~(px_14_6 & be_s1_14);
  assign be_x_14_6 = ~(px_14_7 & be_s1_14);
  assign be_x_14_7 = ~(px_14_8 & be_s1_14);
  assign be_x_14_8 = ~(px_14_9 & be_s1_14);
  assign be_x_14_9 = ~(px_14_10 & be_s1_14);
  assign be_x_15_0 = ~(px_15_1 & be_s1_15);
  assign be_x_15_1 = ~(px_15_2 & be_s1_15);
  assign be_x_15_10 = ~(px_15_11 & be_s1_15);
  assign be_x_15_11 = ~(px_15_12 & be_s1_15);
  assign be_x_15_12 = ~(px_15_13 & be_s1_15);
  assign be_x_15_13 = ~(px_15_14 & be_s1_15);
  assign be_x_15_14 = ~(px_15_15 & be_s1_15);
  assign be_x_15_15 = ~(px_15_16 & be_s1_15);
  assign be_x_15_16 = ~(px_15_17 & be_s1_15);
  assign be_x_15_17 = ~(px_15_18 & be_s1_15);
  assign be_x_15_18 = ~(px_15_19 & be_s1_15);
  assign be_x_15_19 = ~(px_15_20 & be_s1_15);
  assign be_x_15_2 = ~(px_15_3 & be_s1_15);
  assign be_x_15_20 = ~(px_15_21 & be_s1_15);
  assign be_x_15_21 = ~(px_15_22 & be_s1_15);
  assign be_x_15_22 = ~(px_15_23 & be_s1_15);
  assign be_x_15_23 = ~(px_15_24 & be_s1_15);
  assign be_x_15_24 = ~(px_15_25 & be_s1_15);
  assign be_x_15_25 = ~(px_15_26 & be_s1_15);
  assign be_x_15_26 = ~(px_15_27 & be_s1_15);
  assign be_x_15_27 = ~(px_15_28 & be_s1_15);
  assign be_x_15_28 = ~(px_15_29 & be_s1_15);
  assign be_x_15_29 = ~(px_15_30 & be_s1_15);
  assign be_x_15_3 = ~(px_15_4 & be_s1_15);
  assign be_x_15_30 = ~(px_15_31 & be_s1_15);
  assign be_x_15_31 = ~(px_15_32 & be_s1_15);
  assign be_x_15_32 = ~(px_15_33 & be_s1_15);
  assign be_x_15_33 = ~(px_15_34 & be_s1_15);
  assign be_x_15_4 = ~(px_15_5 & be_s1_15);
  assign be_x_15_5 = ~(px_15_6 & be_s1_15);
  assign be_x_15_6 = ~(px_15_7 & be_s1_15);
  assign be_x_15_7 = ~(px_15_8 & be_s1_15);
  assign be_x_15_8 = ~(px_15_9 & be_s1_15);
  assign be_x_15_9 = ~(px_15_10 & be_s1_15);
  assign be_x_16_0 = ~(px_16_1 & be_s1_16);
  assign be_x_16_1 = ~(px_16_2 & be_s1_16);
  assign be_x_16_10 = ~(px_16_11 & be_s1_16);
  assign be_x_16_11 = ~(px_16_12 & be_s1_16);
  assign be_x_16_12 = ~(px_16_13 & be_s1_16);
  assign be_x_16_13 = ~(px_16_14 & be_s1_16);
  assign be_x_16_14 = ~(px_16_15 & be_s1_16);
  assign be_x_16_15 = ~(px_16_16 & be_s1_16);
  assign be_x_16_16 = ~(px_16_17 & be_s1_16);
  assign be_x_16_17 = ~(px_16_18 & be_s1_16);
  assign be_x_16_18 = ~(px_16_19 & be_s1_16);
  assign be_x_16_19 = ~(px_16_20 & be_s1_16);
  assign be_x_16_2 = ~(px_16_3 & be_s1_16);
  assign be_x_16_20 = ~(px_16_21 & be_s1_16);
  assign be_x_16_21 = ~(px_16_22 & be_s1_16);
  assign be_x_16_22 = ~(px_16_23 & be_s1_16);
  assign be_x_16_23 = ~(px_16_24 & be_s1_16);
  assign be_x_16_24 = ~(px_16_25 & be_s1_16);
  assign be_x_16_25 = ~(px_16_26 & be_s1_16);
  assign be_x_16_26 = ~(px_16_27 & be_s1_16);
  assign be_x_16_27 = ~(px_16_28 & be_s1_16);
  assign be_x_16_28 = ~(px_16_29 & be_s1_16);
  assign be_x_16_29 = ~(px_16_30 & be_s1_16);
  assign be_x_16_3 = ~(px_16_4 & be_s1_16);
  assign be_x_16_30 = ~(px_16_31 & be_s1_16);
  assign be_x_16_31 = ~(px_16_32 & be_s1_16);
  assign be_x_16_4 = ~(px_16_5 & be_s1_16);
  assign be_x_16_5 = ~(px_16_6 & be_s1_16);
  assign be_x_16_6 = ~(px_16_7 & be_s1_16);
  assign be_x_16_7 = ~(px_16_8 & be_s1_16);
  assign be_x_16_8 = ~(px_16_9 & be_s1_16);
  assign be_x_16_9 = ~(px_16_10 & be_s1_16);
  assign be_x_1_0 = ~(px_1_1 & be_s1_1);
  assign be_x_1_1 = ~(px_1_2 & be_s1_1);
  assign be_x_1_10 = ~(px_1_11 & be_s1_1);
  assign be_x_1_11 = ~(px_1_12 & be_s1_1);
  assign be_x_1_12 = ~(px_1_13 & be_s1_1);
  assign be_x_1_13 = ~(px_1_14 & be_s1_1);
  assign be_x_1_14 = ~(px_1_15 & be_s1_1);
  assign be_x_1_15 = ~(px_1_16 & be_s1_1);
  assign be_x_1_16 = ~(px_1_17 & be_s1_1);
  assign be_x_1_17 = ~(px_1_18 & be_s1_1);
  assign be_x_1_18 = ~(px_1_19 & be_s1_1);
  assign be_x_1_19 = ~(px_1_20 & be_s1_1);
  assign be_x_1_2 = ~(px_1_3 & be_s1_1);
  assign be_x_1_20 = ~(px_1_21 & be_s1_1);
  assign be_x_1_21 = ~(px_1_22 & be_s1_1);
  assign be_x_1_22 = ~(px_1_23 & be_s1_1);
  assign be_x_1_23 = ~(px_1_24 & be_s1_1);
  assign be_x_1_24 = ~(px_1_25 & be_s1_1);
  assign be_x_1_25 = ~(px_1_26 & be_s1_1);
  assign be_x_1_26 = ~(px_1_27 & be_s1_1);
  assign be_x_1_27 = ~(px_1_28 & be_s1_1);
  assign be_x_1_28 = ~(px_1_29 & be_s1_1);
  assign be_x_1_29 = ~(px_1_30 & be_s1_1);
  assign be_x_1_3 = ~(px_1_4 & be_s1_1);
  assign be_x_1_30 = ~(px_1_31 & be_s1_1);
  assign be_x_1_31 = ~(px_1_32 & be_s1_1);
  assign be_x_1_32 = ~(px_1_33 & be_s1_1);
  assign be_x_1_33 = ~(px_1_34 & be_s1_1);
  assign be_x_1_4 = ~(px_1_5 & be_s1_1);
  assign be_x_1_5 = ~(px_1_6 & be_s1_1);
  assign be_x_1_6 = ~(px_1_7 & be_s1_1);
  assign be_x_1_7 = ~(px_1_8 & be_s1_1);
  assign be_x_1_8 = ~(px_1_9 & be_s1_1);
  assign be_x_1_9 = ~(px_1_10 & be_s1_1);
  assign be_x_2_0 = ~(px_2_1 & be_s1_2);
  assign be_x_2_1 = ~(px_2_2 & be_s1_2);
  assign be_x_2_10 = ~(px_2_11 & be_s1_2);
  assign be_x_2_11 = ~(px_2_12 & be_s1_2);
  assign be_x_2_12 = ~(px_2_13 & be_s1_2);
  assign be_x_2_13 = ~(px_2_14 & be_s1_2);
  assign be_x_2_14 = ~(px_2_15 & be_s1_2);
  assign be_x_2_15 = ~(px_2_16 & be_s1_2);
  assign be_x_2_16 = ~(px_2_17 & be_s1_2);
  assign be_x_2_17 = ~(px_2_18 & be_s1_2);
  assign be_x_2_18 = ~(px_2_19 & be_s1_2);
  assign be_x_2_19 = ~(px_2_20 & be_s1_2);
  assign be_x_2_2 = ~(px_2_3 & be_s1_2);
  assign be_x_2_20 = ~(px_2_21 & be_s1_2);
  assign be_x_2_21 = ~(px_2_22 & be_s1_2);
  assign be_x_2_22 = ~(px_2_23 & be_s1_2);
  assign be_x_2_23 = ~(px_2_24 & be_s1_2);
  assign be_x_2_24 = ~(px_2_25 & be_s1_2);
  assign be_x_2_25 = ~(px_2_26 & be_s1_2);
  assign be_x_2_26 = ~(px_2_27 & be_s1_2);
  assign be_x_2_27 = ~(px_2_28 & be_s1_2);
  assign be_x_2_28 = ~(px_2_29 & be_s1_2);
  assign be_x_2_29 = ~(px_2_30 & be_s1_2);
  assign be_x_2_3 = ~(px_2_4 & be_s1_2);
  assign be_x_2_30 = ~(px_2_31 & be_s1_2);
  assign be_x_2_31 = ~(px_2_32 & be_s1_2);
  assign be_x_2_32 = ~(px_2_33 & be_s1_2);
  assign be_x_2_33 = ~(px_2_34 & be_s1_2);
  assign be_x_2_4 = ~(px_2_5 & be_s1_2);
  assign be_x_2_5 = ~(px_2_6 & be_s1_2);
  assign be_x_2_6 = ~(px_2_7 & be_s1_2);
  assign be_x_2_7 = ~(px_2_8 & be_s1_2);
  assign be_x_2_8 = ~(px_2_9 & be_s1_2);
  assign be_x_2_9 = ~(px_2_10 & be_s1_2);
  assign be_x_3_0 = ~(px_3_1 & be_s1_3);
  assign be_x_3_1 = ~(px_3_2 & be_s1_3);
  assign be_x_3_10 = ~(px_3_11 & be_s1_3);
  assign be_x_3_11 = ~(px_3_12 & be_s1_3);
  assign be_x_3_12 = ~(px_3_13 & be_s1_3);
  assign be_x_3_13 = ~(px_3_14 & be_s1_3);
  assign be_x_3_14 = ~(px_3_15 & be_s1_3);
  assign be_x_3_15 = ~(px_3_16 & be_s1_3);
  assign be_x_3_16 = ~(px_3_17 & be_s1_3);
  assign be_x_3_17 = ~(px_3_18 & be_s1_3);
  assign be_x_3_18 = ~(px_3_19 & be_s1_3);
  assign be_x_3_19 = ~(px_3_20 & be_s1_3);
  assign be_x_3_2 = ~(px_3_3 & be_s1_3);
  assign be_x_3_20 = ~(px_3_21 & be_s1_3);
  assign be_x_3_21 = ~(px_3_22 & be_s1_3);
  assign be_x_3_22 = ~(px_3_23 & be_s1_3);
  assign be_x_3_23 = ~(px_3_24 & be_s1_3);
  assign be_x_3_24 = ~(px_3_25 & be_s1_3);
  assign be_x_3_25 = ~(px_3_26 & be_s1_3);
  assign be_x_3_26 = ~(px_3_27 & be_s1_3);
  assign be_x_3_27 = ~(px_3_28 & be_s1_3);
  assign be_x_3_28 = ~(px_3_29 & be_s1_3);
  assign be_x_3_29 = ~(px_3_30 & be_s1_3);
  assign be_x_3_3 = ~(px_3_4 & be_s1_3);
  assign be_x_3_30 = ~(px_3_31 & be_s1_3);
  assign be_x_3_31 = ~(px_3_32 & be_s1_3);
  assign be_x_3_32 = ~(px_3_33 & be_s1_3);
  assign be_x_3_33 = ~(px_3_34 & be_s1_3);
  assign be_x_3_4 = ~(px_3_5 & be_s1_3);
  assign be_x_3_5 = ~(px_3_6 & be_s1_3);
  assign be_x_3_6 = ~(px_3_7 & be_s1_3);
  assign be_x_3_7 = ~(px_3_8 & be_s1_3);
  assign be_x_3_8 = ~(px_3_9 & be_s1_3);
  assign be_x_3_9 = ~(px_3_10 & be_s1_3);
  assign be_x_4_0 = ~(px_4_1 & be_s1_4);
  assign be_x_4_1 = ~(px_4_2 & be_s1_4);
  assign be_x_4_10 = ~(px_4_11 & be_s1_4);
  assign be_x_4_11 = ~(px_4_12 & be_s1_4);
  assign be_x_4_12 = ~(px_4_13 & be_s1_4);
  assign be_x_4_13 = ~(px_4_14 & be_s1_4);
  assign be_x_4_14 = ~(px_4_15 & be_s1_4);
  assign be_x_4_15 = ~(px_4_16 & be_s1_4);
  assign be_x_4_16 = ~(px_4_17 & be_s1_4);
  assign be_x_4_17 = ~(px_4_18 & be_s1_4);
  assign be_x_4_18 = ~(px_4_19 & be_s1_4);
  assign be_x_4_19 = ~(px_4_20 & be_s1_4);
  assign be_x_4_2 = ~(px_4_3 & be_s1_4);
  assign be_x_4_20 = ~(px_4_21 & be_s1_4);
  assign be_x_4_21 = ~(px_4_22 & be_s1_4);
  assign be_x_4_22 = ~(px_4_23 & be_s1_4);
  assign be_x_4_23 = ~(px_4_24 & be_s1_4);
  assign be_x_4_24 = ~(px_4_25 & be_s1_4);
  assign be_x_4_25 = ~(px_4_26 & be_s1_4);
  assign be_x_4_26 = ~(px_4_27 & be_s1_4);
  assign be_x_4_27 = ~(px_4_28 & be_s1_4);
  assign be_x_4_28 = ~(px_4_29 & be_s1_4);
  assign be_x_4_29 = ~(px_4_30 & be_s1_4);
  assign be_x_4_3 = ~(px_4_4 & be_s1_4);
  assign be_x_4_30 = ~(px_4_31 & be_s1_4);
  assign be_x_4_31 = ~(px_4_32 & be_s1_4);
  assign be_x_4_32 = ~(px_4_33 & be_s1_4);
  assign be_x_4_33 = ~(px_4_34 & be_s1_4);
  assign be_x_4_4 = ~(px_4_5 & be_s1_4);
  assign be_x_4_5 = ~(px_4_6 & be_s1_4);
  assign be_x_4_6 = ~(px_4_7 & be_s1_4);
  assign be_x_4_7 = ~(px_4_8 & be_s1_4);
  assign be_x_4_8 = ~(px_4_9 & be_s1_4);
  assign be_x_4_9 = ~(px_4_10 & be_s1_4);
  assign be_x_5_0 = ~(px_5_1 & be_s1_5);
  assign be_x_5_1 = ~(px_5_2 & be_s1_5);
  assign be_x_5_10 = ~(px_5_11 & be_s1_5);
  assign be_x_5_11 = ~(px_5_12 & be_s1_5);
  assign be_x_5_12 = ~(px_5_13 & be_s1_5);
  assign be_x_5_13 = ~(px_5_14 & be_s1_5);
  assign be_x_5_14 = ~(px_5_15 & be_s1_5);
  assign be_x_5_15 = ~(px_5_16 & be_s1_5);
  assign be_x_5_16 = ~(px_5_17 & be_s1_5);
  assign be_x_5_17 = ~(px_5_18 & be_s1_5);
  assign be_x_5_18 = ~(px_5_19 & be_s1_5);
  assign be_x_5_19 = ~(px_5_20 & be_s1_5);
  assign be_x_5_2 = ~(px_5_3 & be_s1_5);
  assign be_x_5_20 = ~(px_5_21 & be_s1_5);
  assign be_x_5_21 = ~(px_5_22 & be_s1_5);
  assign be_x_5_22 = ~(px_5_23 & be_s1_5);
  assign be_x_5_23 = ~(px_5_24 & be_s1_5);
  assign be_x_5_24 = ~(px_5_25 & be_s1_5);
  assign be_x_5_25 = ~(px_5_26 & be_s1_5);
  assign be_x_5_26 = ~(px_5_27 & be_s1_5);
  assign be_x_5_27 = ~(px_5_28 & be_s1_5);
  assign be_x_5_28 = ~(px_5_29 & be_s1_5);
  assign be_x_5_29 = ~(px_5_30 & be_s1_5);
  assign be_x_5_3 = ~(px_5_4 & be_s1_5);
  assign be_x_5_30 = ~(px_5_31 & be_s1_5);
  assign be_x_5_31 = ~(px_5_32 & be_s1_5);
  assign be_x_5_32 = ~(px_5_33 & be_s1_5);
  assign be_x_5_33 = ~(px_5_34 & be_s1_5);
  assign be_x_5_4 = ~(px_5_5 & be_s1_5);
  assign be_x_5_5 = ~(px_5_6 & be_s1_5);
  assign be_x_5_6 = ~(px_5_7 & be_s1_5);
  assign be_x_5_7 = ~(px_5_8 & be_s1_5);
  assign be_x_5_8 = ~(px_5_9 & be_s1_5);
  assign be_x_5_9 = ~(px_5_10 & be_s1_5);
  assign be_x_6_0 = ~(px_6_1 & be_s1_6);
  assign be_x_6_1 = ~(px_6_2 & be_s1_6);
  assign be_x_6_10 = ~(px_6_11 & be_s1_6);
  assign be_x_6_11 = ~(px_6_12 & be_s1_6);
  assign be_x_6_12 = ~(px_6_13 & be_s1_6);
  assign be_x_6_13 = ~(px_6_14 & be_s1_6);
  assign be_x_6_14 = ~(px_6_15 & be_s1_6);
  assign be_x_6_15 = ~(px_6_16 & be_s1_6);
  assign be_x_6_16 = ~(px_6_17 & be_s1_6);
  assign be_x_6_17 = ~(px_6_18 & be_s1_6);
  assign be_x_6_18 = ~(px_6_19 & be_s1_6);
  assign be_x_6_19 = ~(px_6_20 & be_s1_6);
  assign be_x_6_2 = ~(px_6_3 & be_s1_6);
  assign be_x_6_20 = ~(px_6_21 & be_s1_6);
  assign be_x_6_21 = ~(px_6_22 & be_s1_6);
  assign be_x_6_22 = ~(px_6_23 & be_s1_6);
  assign be_x_6_23 = ~(px_6_24 & be_s1_6);
  assign be_x_6_24 = ~(px_6_25 & be_s1_6);
  assign be_x_6_25 = ~(px_6_26 & be_s1_6);
  assign be_x_6_26 = ~(px_6_27 & be_s1_6);
  assign be_x_6_27 = ~(px_6_28 & be_s1_6);
  assign be_x_6_28 = ~(px_6_29 & be_s1_6);
  assign be_x_6_29 = ~(px_6_30 & be_s1_6);
  assign be_x_6_3 = ~(px_6_4 & be_s1_6);
  assign be_x_6_30 = ~(px_6_31 & be_s1_6);
  assign be_x_6_31 = ~(px_6_32 & be_s1_6);
  assign be_x_6_32 = ~(px_6_33 & be_s1_6);
  assign be_x_6_33 = ~(px_6_34 & be_s1_6);
  assign be_x_6_4 = ~(px_6_5 & be_s1_6);
  assign be_x_6_5 = ~(px_6_6 & be_s1_6);
  assign be_x_6_6 = ~(px_6_7 & be_s1_6);
  assign be_x_6_7 = ~(px_6_8 & be_s1_6);
  assign be_x_6_8 = ~(px_6_9 & be_s1_6);
  assign be_x_6_9 = ~(px_6_10 & be_s1_6);
  assign be_x_7_0 = ~(px_7_1 & be_s1_7);
  assign be_x_7_1 = ~(px_7_2 & be_s1_7);
  assign be_x_7_10 = ~(px_7_11 & be_s1_7);
  assign be_x_7_11 = ~(px_7_12 & be_s1_7);
  assign be_x_7_12 = ~(px_7_13 & be_s1_7);
  assign be_x_7_13 = ~(px_7_14 & be_s1_7);
  assign be_x_7_14 = ~(px_7_15 & be_s1_7);
  assign be_x_7_15 = ~(px_7_16 & be_s1_7);
  assign be_x_7_16 = ~(px_7_17 & be_s1_7);
  assign be_x_7_17 = ~(px_7_18 & be_s1_7);
  assign be_x_7_18 = ~(px_7_19 & be_s1_7);
  assign be_x_7_19 = ~(px_7_20 & be_s1_7);
  assign be_x_7_2 = ~(px_7_3 & be_s1_7);
  assign be_x_7_20 = ~(px_7_21 & be_s1_7);
  assign be_x_7_21 = ~(px_7_22 & be_s1_7);
  assign be_x_7_22 = ~(px_7_23 & be_s1_7);
  assign be_x_7_23 = ~(px_7_24 & be_s1_7);
  assign be_x_7_24 = ~(px_7_25 & be_s1_7);
  assign be_x_7_25 = ~(px_7_26 & be_s1_7);
  assign be_x_7_26 = ~(px_7_27 & be_s1_7);
  assign be_x_7_27 = ~(px_7_28 & be_s1_7);
  assign be_x_7_28 = ~(px_7_29 & be_s1_7);
  assign be_x_7_29 = ~(px_7_30 & be_s1_7);
  assign be_x_7_3 = ~(px_7_4 & be_s1_7);
  assign be_x_7_30 = ~(px_7_31 & be_s1_7);
  assign be_x_7_31 = ~(px_7_32 & be_s1_7);
  assign be_x_7_32 = ~(px_7_33 & be_s1_7);
  assign be_x_7_33 = ~(px_7_34 & be_s1_7);
  assign be_x_7_4 = ~(px_7_5 & be_s1_7);
  assign be_x_7_5 = ~(px_7_6 & be_s1_7);
  assign be_x_7_6 = ~(px_7_7 & be_s1_7);
  assign be_x_7_7 = ~(px_7_8 & be_s1_7);
  assign be_x_7_8 = ~(px_7_9 & be_s1_7);
  assign be_x_7_9 = ~(px_7_10 & be_s1_7);
  assign be_x_8_0 = ~(px_8_1 & be_s1_8);
  assign be_x_8_1 = ~(px_8_2 & be_s1_8);
  assign be_x_8_10 = ~(px_8_11 & be_s1_8);
  assign be_x_8_11 = ~(px_8_12 & be_s1_8);
  assign be_x_8_12 = ~(px_8_13 & be_s1_8);
  assign be_x_8_13 = ~(px_8_14 & be_s1_8);
  assign be_x_8_14 = ~(px_8_15 & be_s1_8);
  assign be_x_8_15 = ~(px_8_16 & be_s1_8);
  assign be_x_8_16 = ~(px_8_17 & be_s1_8);
  assign be_x_8_17 = ~(px_8_18 & be_s1_8);
  assign be_x_8_18 = ~(px_8_19 & be_s1_8);
  assign be_x_8_19 = ~(px_8_20 & be_s1_8);
  assign be_x_8_2 = ~(px_8_3 & be_s1_8);
  assign be_x_8_20 = ~(px_8_21 & be_s1_8);
  assign be_x_8_21 = ~(px_8_22 & be_s1_8);
  assign be_x_8_22 = ~(px_8_23 & be_s1_8);
  assign be_x_8_23 = ~(px_8_24 & be_s1_8);
  assign be_x_8_24 = ~(px_8_25 & be_s1_8);
  assign be_x_8_25 = ~(px_8_26 & be_s1_8);
  assign be_x_8_26 = ~(px_8_27 & be_s1_8);
  assign be_x_8_27 = ~(px_8_28 & be_s1_8);
  assign be_x_8_28 = ~(px_8_29 & be_s1_8);
  assign be_x_8_29 = ~(px_8_30 & be_s1_8);
  assign be_x_8_3 = ~(px_8_4 & be_s1_8);
  assign be_x_8_30 = ~(px_8_31 & be_s1_8);
  assign be_x_8_31 = ~(px_8_32 & be_s1_8);
  assign be_x_8_32 = ~(px_8_33 & be_s1_8);
  assign be_x_8_33 = ~(px_8_34 & be_s1_8);
  assign be_x_8_4 = ~(px_8_5 & be_s1_8);
  assign be_x_8_5 = ~(px_8_6 & be_s1_8);
  assign be_x_8_6 = ~(px_8_7 & be_s1_8);
  assign be_x_8_7 = ~(px_8_8 & be_s1_8);
  assign be_x_8_8 = ~(px_8_9 & be_s1_8);
  assign be_x_8_9 = ~(px_8_10 & be_s1_8);
  assign be_x_9_0 = ~(px_9_1 & be_s1_9);
  assign be_x_9_1 = ~(px_9_2 & be_s1_9);
  assign be_x_9_10 = ~(px_9_11 & be_s1_9);
  assign be_x_9_11 = ~(px_9_12 & be_s1_9);
  assign be_x_9_12 = ~(px_9_13 & be_s1_9);
  assign be_x_9_13 = ~(px_9_14 & be_s1_9);
  assign be_x_9_14 = ~(px_9_15 & be_s1_9);
  assign be_x_9_15 = ~(px_9_16 & be_s1_9);
  assign be_x_9_16 = ~(px_9_17 & be_s1_9);
  assign be_x_9_17 = ~(px_9_18 & be_s1_9);
  assign be_x_9_18 = ~(px_9_19 & be_s1_9);
  assign be_x_9_19 = ~(px_9_20 & be_s1_9);
  assign be_x_9_2 = ~(px_9_3 & be_s1_9);
  assign be_x_9_20 = ~(px_9_21 & be_s1_9);
  assign be_x_9_21 = ~(px_9_22 & be_s1_9);
  assign be_x_9_22 = ~(px_9_23 & be_s1_9);
  assign be_x_9_23 = ~(px_9_24 & be_s1_9);
  assign be_x_9_24 = ~(px_9_25 & be_s1_9);
  assign be_x_9_25 = ~(px_9_26 & be_s1_9);
  assign be_x_9_26 = ~(px_9_27 & be_s1_9);
  assign be_x_9_27 = ~(px_9_28 & be_s1_9);
  assign be_x_9_28 = ~(px_9_29 & be_s1_9);
  assign be_x_9_29 = ~(px_9_30 & be_s1_9);
  assign be_x_9_3 = ~(px_9_4 & be_s1_9);
  assign be_x_9_30 = ~(px_9_31 & be_s1_9);
  assign be_x_9_31 = ~(px_9_32 & be_s1_9);
  assign be_x_9_32 = ~(px_9_33 & be_s1_9);
  assign be_x_9_33 = ~(px_9_34 & be_s1_9);
  assign be_x_9_4 = ~(px_9_5 & be_s1_9);
  assign be_x_9_5 = ~(px_9_6 & be_s1_9);
  assign be_x_9_6 = ~(px_9_7 & be_s1_9);
  assign be_x_9_7 = ~(px_9_8 & be_s1_9);
  assign be_x_9_8 = ~(px_9_9 & be_s1_9);
  assign be_x_9_9 = ~(px_9_10 & be_s1_9);
  assign not_pp_0_35 = ~pp_0_33;
  assign not_pp_10_53 = ~pp_10_53;
  assign not_pp_11_55 = ~pp_11_55;
  assign not_pp_12_57 = ~pp_12_57;
  assign not_pp_13_59 = ~pp_13_59;
  assign not_pp_14_61 = ~pp_14_61;
  assign not_pp_15_63 = ~pp_15_63;
  assign not_pp_1_35 = ~pp_1_35;
  assign not_pp_2_37 = ~pp_2_37;
  assign not_pp_3_39 = ~pp_3_39;
  assign not_pp_4_41 = ~pp_4_41;
  assign not_pp_5_43 = ~pp_5_43;
  assign not_pp_6_45 = ~pp_6_45;
  assign not_pp_7_47 = ~pp_7_47;
  assign not_pp_8_49 = ~pp_8_49;
  assign not_pp_9_51 = ~pp_9_51;
  assign ny_0 = ~multiplier[0];
  assign ny_1 = ~multiplier[1];
  assign ny_10 = ~multiplier[10];
  assign ny_11 = ~multiplier[11];
  assign ny_12 = ~multiplier[12];
  assign ny_13 = ~multiplier[13];
  assign ny_14 = ~multiplier[14];
  assign ny_15 = ~multiplier[15];
  assign ny_16 = ~multiplier[16];
  assign ny_17 = ~multiplier[17];
  assign ny_18 = ~multiplier[18];
  assign ny_19 = ~multiplier[19];
  assign ny_2 = ~multiplier[2];
  assign ny_20 = ~multiplier[20];
  assign ny_21 = ~multiplier[21];
  assign ny_22 = ~multiplier[22];
  assign ny_23 = ~multiplier[23];
  assign ny_24 = ~multiplier[24];
  assign ny_25 = ~multiplier[25];
  assign ny_26 = ~multiplier[26];
  assign ny_27 = ~multiplier[27];
  assign ny_28 = ~multiplier[28];
  assign ny_29 = ~multiplier[29];
  assign ny_3 = ~multiplier[3];
  assign ny_30 = ~multiplier[30];
  assign ny_31 = ~multiplier[31];
  assign ny_4 = ~multiplier[4];
  assign ny_5 = ~multiplier[5];
  assign ny_6 = ~multiplier[6];
  assign ny_7 = ~multiplier[7];
  assign ny_8 = ~multiplier[8];
  assign ny_9 = ~multiplier[9];
  assign one = 1'b1;
  assign pp_0_0 = ~(be_2x_0_0 & be_x_0_0);
  assign pp_0_1 = ~(be_2x_0_1 & be_x_0_1);
  assign pp_0_10 = ~(be_2x_0_10 & be_x_0_10);
  assign pp_0_11 = ~(be_2x_0_11 & be_x_0_11);
  assign pp_0_12 = ~(be_2x_0_12 & be_x_0_12);
  assign pp_0_13 = ~(be_2x_0_13 & be_x_0_13);
  assign pp_0_14 = ~(be_2x_0_14 & be_x_0_14);
  assign pp_0_15 = ~(be_2x_0_15 & be_x_0_15);
  assign pp_0_16 = ~(be_2x_0_16 & be_x_0_16);
  assign pp_0_17 = ~(be_2x_0_17 & be_x_0_17);
  assign pp_0_18 = ~(be_2x_0_18 & be_x_0_18);
  assign pp_0_19 = ~(be_2x_0_19 & be_x_0_19);
  assign pp_0_2 = ~(be_2x_0_2 & be_x_0_2);
  assign pp_0_20 = ~(be_2x_0_20 & be_x_0_20);
  assign pp_0_21 = ~(be_2x_0_21 & be_x_0_21);
  assign pp_0_22 = ~(be_2x_0_22 & be_x_0_22);
  assign pp_0_23 = ~(be_2x_0_23 & be_x_0_23);
  assign pp_0_24 = ~(be_2x_0_24 & be_x_0_24);
  assign pp_0_25 = ~(be_2x_0_25 & be_x_0_25);
  assign pp_0_26 = ~(be_2x_0_26 & be_x_0_26);
  assign pp_0_27 = ~(be_2x_0_27 & be_x_0_27);
  assign pp_0_28 = ~(be_2x_0_28 & be_x_0_28);
  assign pp_0_29 = ~(be_2x_0_29 & be_x_0_29);
  assign pp_0_3 = ~(be_2x_0_3 & be_x_0_3);
  assign pp_0_30 = ~(be_2x_0_30 & be_x_0_30);
  assign pp_0_31 = ~(be_2x_0_31 & be_x_0_31);
  assign pp_0_32 = ~(be_2x_0_32 & be_x_0_32);
  assign pp_0_33 = ~(be_2x_0_33 & be_x_0_33);
  assign pp_0_4 = ~(be_2x_0_4 & be_x_0_4);
  assign pp_0_5 = ~(be_2x_0_5 & be_x_0_5);
  assign pp_0_6 = ~(be_2x_0_6 & be_x_0_6);
  assign pp_0_7 = ~(be_2x_0_7 & be_x_0_7);
  assign pp_0_8 = ~(be_2x_0_8 & be_x_0_8);
  assign pp_0_9 = ~(be_2x_0_9 & be_x_0_9);
  assign pp_10_20 = ~(be_2x_10_0 & be_x_10_0);
  assign pp_10_21 = ~(be_2x_10_1 & be_x_10_1);
  assign pp_10_22 = ~(be_2x_10_2 & be_x_10_2);
  assign pp_10_23 = ~(be_2x_10_3 & be_x_10_3);
  assign pp_10_24 = ~(be_2x_10_4 & be_x_10_4);
  assign pp_10_25 = ~(be_2x_10_5 & be_x_10_5);
  assign pp_10_26 = ~(be_2x_10_6 & be_x_10_6);
  assign pp_10_27 = ~(be_2x_10_7 & be_x_10_7);
  assign pp_10_28 = ~(be_2x_10_8 & be_x_10_8);
  assign pp_10_29 = ~(be_2x_10_9 & be_x_10_9);
  assign pp_10_30 = ~(be_2x_10_10 & be_x_10_10);
  assign pp_10_31 = ~(be_2x_10_11 & be_x_10_11);
  assign pp_10_32 = ~(be_2x_10_12 & be_x_10_12);
  assign pp_10_33 = ~(be_2x_10_13 & be_x_10_13);
  assign pp_10_34 = ~(be_2x_10_14 & be_x_10_14);
  assign pp_10_35 = ~(be_2x_10_15 & be_x_10_15);
  assign pp_10_36 = ~(be_2x_10_16 & be_x_10_16);
  assign pp_10_37 = ~(be_2x_10_17 & be_x_10_17);
  assign pp_10_38 = ~(be_2x_10_18 & be_x_10_18);
  assign pp_10_39 = ~(be_2x_10_19 & be_x_10_19);
  assign pp_10_40 = ~(be_2x_10_20 & be_x_10_20);
  assign pp_10_41 = ~(be_2x_10_21 & be_x_10_21);
  assign pp_10_42 = ~(be_2x_10_22 & be_x_10_22);
  assign pp_10_43 = ~(be_2x_10_23 & be_x_10_23);
  assign pp_10_44 = ~(be_2x_10_24 & be_x_10_24);
  assign pp_10_45 = ~(be_2x_10_25 & be_x_10_25);
  assign pp_10_46 = ~(be_2x_10_26 & be_x_10_26);
  assign pp_10_47 = ~(be_2x_10_27 & be_x_10_27);
  assign pp_10_48 = ~(be_2x_10_28 & be_x_10_28);
  assign pp_10_49 = ~(be_2x_10_29 & be_x_10_29);
  assign pp_10_50 = ~(be_2x_10_30 & be_x_10_30);
  assign pp_10_51 = ~(be_2x_10_31 & be_x_10_31);
  assign pp_10_52 = ~(be_2x_10_32 & be_x_10_32);
  assign pp_10_53 = ~(be_2x_10_33 & be_x_10_33);
  assign pp_11_22 = ~(be_2x_11_0 & be_x_11_0);
  assign pp_11_23 = ~(be_2x_11_1 & be_x_11_1);
  assign pp_11_24 = ~(be_2x_11_2 & be_x_11_2);
  assign pp_11_25 = ~(be_2x_11_3 & be_x_11_3);
  assign pp_11_26 = ~(be_2x_11_4 & be_x_11_4);
  assign pp_11_27 = ~(be_2x_11_5 & be_x_11_5);
  assign pp_11_28 = ~(be_2x_11_6 & be_x_11_6);
  assign pp_11_29 = ~(be_2x_11_7 & be_x_11_7);
  assign pp_11_30 = ~(be_2x_11_8 & be_x_11_8);
  assign pp_11_31 = ~(be_2x_11_9 & be_x_11_9);
  assign pp_11_32 = ~(be_2x_11_10 & be_x_11_10);
  assign pp_11_33 = ~(be_2x_11_11 & be_x_11_11);
  assign pp_11_34 = ~(be_2x_11_12 & be_x_11_12);
  assign pp_11_35 = ~(be_2x_11_13 & be_x_11_13);
  assign pp_11_36 = ~(be_2x_11_14 & be_x_11_14);
  assign pp_11_37 = ~(be_2x_11_15 & be_x_11_15);
  assign pp_11_38 = ~(be_2x_11_16 & be_x_11_16);
  assign pp_11_39 = ~(be_2x_11_17 & be_x_11_17);
  assign pp_11_40 = ~(be_2x_11_18 & be_x_11_18);
  assign pp_11_41 = ~(be_2x_11_19 & be_x_11_19);
  assign pp_11_42 = ~(be_2x_11_20 & be_x_11_20);
  assign pp_11_43 = ~(be_2x_11_21 & be_x_11_21);
  assign pp_11_44 = ~(be_2x_11_22 & be_x_11_22);
  assign pp_11_45 = ~(be_2x_11_23 & be_x_11_23);
  assign pp_11_46 = ~(be_2x_11_24 & be_x_11_24);
  assign pp_11_47 = ~(be_2x_11_25 & be_x_11_25);
  assign pp_11_48 = ~(be_2x_11_26 & be_x_11_26);
  assign pp_11_49 = ~(be_2x_11_27 & be_x_11_27);
  assign pp_11_50 = ~(be_2x_11_28 & be_x_11_28);
  assign pp_11_51 = ~(be_2x_11_29 & be_x_11_29);
  assign pp_11_52 = ~(be_2x_11_30 & be_x_11_30);
  assign pp_11_53 = ~(be_2x_11_31 & be_x_11_31);
  assign pp_11_54 = ~(be_2x_11_32 & be_x_11_32);
  assign pp_11_55 = ~(be_2x_11_33 & be_x_11_33);
  assign pp_12_24 = ~(be_2x_12_0 & be_x_12_0);
  assign pp_12_25 = ~(be_2x_12_1 & be_x_12_1);
  assign pp_12_26 = ~(be_2x_12_2 & be_x_12_2);
  assign pp_12_27 = ~(be_2x_12_3 & be_x_12_3);
  assign pp_12_28 = ~(be_2x_12_4 & be_x_12_4);
  assign pp_12_29 = ~(be_2x_12_5 & be_x_12_5);
  assign pp_12_30 = ~(be_2x_12_6 & be_x_12_6);
  assign pp_12_31 = ~(be_2x_12_7 & be_x_12_7);
  assign pp_12_32 = ~(be_2x_12_8 & be_x_12_8);
  assign pp_12_33 = ~(be_2x_12_9 & be_x_12_9);
  assign pp_12_34 = ~(be_2x_12_10 & be_x_12_10);
  assign pp_12_35 = ~(be_2x_12_11 & be_x_12_11);
  assign pp_12_36 = ~(be_2x_12_12 & be_x_12_12);
  assign pp_12_37 = ~(be_2x_12_13 & be_x_12_13);
  assign pp_12_38 = ~(be_2x_12_14 & be_x_12_14);
  assign pp_12_39 = ~(be_2x_12_15 & be_x_12_15);
  assign pp_12_40 = ~(be_2x_12_16 & be_x_12_16);
  assign pp_12_41 = ~(be_2x_12_17 & be_x_12_17);
  assign pp_12_42 = ~(be_2x_12_18 & be_x_12_18);
  assign pp_12_43 = ~(be_2x_12_19 & be_x_12_19);
  assign pp_12_44 = ~(be_2x_12_20 & be_x_12_20);
  assign pp_12_45 = ~(be_2x_12_21 & be_x_12_21);
  assign pp_12_46 = ~(be_2x_12_22 & be_x_12_22);
  assign pp_12_47 = ~(be_2x_12_23 & be_x_12_23);
  assign pp_12_48 = ~(be_2x_12_24 & be_x_12_24);
  assign pp_12_49 = ~(be_2x_12_25 & be_x_12_25);
  assign pp_12_50 = ~(be_2x_12_26 & be_x_12_26);
  assign pp_12_51 = ~(be_2x_12_27 & be_x_12_27);
  assign pp_12_52 = ~(be_2x_12_28 & be_x_12_28);
  assign pp_12_53 = ~(be_2x_12_29 & be_x_12_29);
  assign pp_12_54 = ~(be_2x_12_30 & be_x_12_30);
  assign pp_12_55 = ~(be_2x_12_31 & be_x_12_31);
  assign pp_12_56 = ~(be_2x_12_32 & be_x_12_32);
  assign pp_12_57 = ~(be_2x_12_33 & be_x_12_33);
  assign pp_13_26 = ~(be_2x_13_0 & be_x_13_0);
  assign pp_13_27 = ~(be_2x_13_1 & be_x_13_1);
  assign pp_13_28 = ~(be_2x_13_2 & be_x_13_2);
  assign pp_13_29 = ~(be_2x_13_3 & be_x_13_3);
  assign pp_13_30 = ~(be_2x_13_4 & be_x_13_4);
  assign pp_13_31 = ~(be_2x_13_5 & be_x_13_5);
  assign pp_13_32 = ~(be_2x_13_6 & be_x_13_6);
  assign pp_13_33 = ~(be_2x_13_7 & be_x_13_7);
  assign pp_13_34 = ~(be_2x_13_8 & be_x_13_8);
  assign pp_13_35 = ~(be_2x_13_9 & be_x_13_9);
  assign pp_13_36 = ~(be_2x_13_10 & be_x_13_10);
  assign pp_13_37 = ~(be_2x_13_11 & be_x_13_11);
  assign pp_13_38 = ~(be_2x_13_12 & be_x_13_12);
  assign pp_13_39 = ~(be_2x_13_13 & be_x_13_13);
  assign pp_13_40 = ~(be_2x_13_14 & be_x_13_14);
  assign pp_13_41 = ~(be_2x_13_15 & be_x_13_15);
  assign pp_13_42 = ~(be_2x_13_16 & be_x_13_16);
  assign pp_13_43 = ~(be_2x_13_17 & be_x_13_17);
  assign pp_13_44 = ~(be_2x_13_18 & be_x_13_18);
  assign pp_13_45 = ~(be_2x_13_19 & be_x_13_19);
  assign pp_13_46 = ~(be_2x_13_20 & be_x_13_20);
  assign pp_13_47 = ~(be_2x_13_21 & be_x_13_21);
  assign pp_13_48 = ~(be_2x_13_22 & be_x_13_22);
  assign pp_13_49 = ~(be_2x_13_23 & be_x_13_23);
  assign pp_13_50 = ~(be_2x_13_24 & be_x_13_24);
  assign pp_13_51 = ~(be_2x_13_25 & be_x_13_25);
  assign pp_13_52 = ~(be_2x_13_26 & be_x_13_26);
  assign pp_13_53 = ~(be_2x_13_27 & be_x_13_27);
  assign pp_13_54 = ~(be_2x_13_28 & be_x_13_28);
  assign pp_13_55 = ~(be_2x_13_29 & be_x_13_29);
  assign pp_13_56 = ~(be_2x_13_30 & be_x_13_30);
  assign pp_13_57 = ~(be_2x_13_31 & be_x_13_31);
  assign pp_13_58 = ~(be_2x_13_32 & be_x_13_32);
  assign pp_13_59 = ~(be_2x_13_33 & be_x_13_33);
  assign pp_14_28 = ~(be_2x_14_0 & be_x_14_0);
  assign pp_14_29 = ~(be_2x_14_1 & be_x_14_1);
  assign pp_14_30 = ~(be_2x_14_2 & be_x_14_2);
  assign pp_14_31 = ~(be_2x_14_3 & be_x_14_3);
  assign pp_14_32 = ~(be_2x_14_4 & be_x_14_4);
  assign pp_14_33 = ~(be_2x_14_5 & be_x_14_5);
  assign pp_14_34 = ~(be_2x_14_6 & be_x_14_6);
  assign pp_14_35 = ~(be_2x_14_7 & be_x_14_7);
  assign pp_14_36 = ~(be_2x_14_8 & be_x_14_8);
  assign pp_14_37 = ~(be_2x_14_9 & be_x_14_9);
  assign pp_14_38 = ~(be_2x_14_10 & be_x_14_10);
  assign pp_14_39 = ~(be_2x_14_11 & be_x_14_11);
  assign pp_14_40 = ~(be_2x_14_12 & be_x_14_12);
  assign pp_14_41 = ~(be_2x_14_13 & be_x_14_13);
  assign pp_14_42 = ~(be_2x_14_14 & be_x_14_14);
  assign pp_14_43 = ~(be_2x_14_15 & be_x_14_15);
  assign pp_14_44 = ~(be_2x_14_16 & be_x_14_16);
  assign pp_14_45 = ~(be_2x_14_17 & be_x_14_17);
  assign pp_14_46 = ~(be_2x_14_18 & be_x_14_18);
  assign pp_14_47 = ~(be_2x_14_19 & be_x_14_19);
  assign pp_14_48 = ~(be_2x_14_20 & be_x_14_20);
  assign pp_14_49 = ~(be_2x_14_21 & be_x_14_21);
  assign pp_14_50 = ~(be_2x_14_22 & be_x_14_22);
  assign pp_14_51 = ~(be_2x_14_23 & be_x_14_23);
  assign pp_14_52 = ~(be_2x_14_24 & be_x_14_24);
  assign pp_14_53 = ~(be_2x_14_25 & be_x_14_25);
  assign pp_14_54 = ~(be_2x_14_26 & be_x_14_26);
  assign pp_14_55 = ~(be_2x_14_27 & be_x_14_27);
  assign pp_14_56 = ~(be_2x_14_28 & be_x_14_28);
  assign pp_14_57 = ~(be_2x_14_29 & be_x_14_29);
  assign pp_14_58 = ~(be_2x_14_30 & be_x_14_30);
  assign pp_14_59 = ~(be_2x_14_31 & be_x_14_31);
  assign pp_14_60 = ~(be_2x_14_32 & be_x_14_32);
  assign pp_14_61 = ~(be_2x_14_33 & be_x_14_33);
  assign pp_15_30 = ~(be_2x_15_0 & be_x_15_0);
  assign pp_15_31 = ~(be_2x_15_1 & be_x_15_1);
  assign pp_15_32 = ~(be_2x_15_2 & be_x_15_2);
  assign pp_15_33 = ~(be_2x_15_3 & be_x_15_3);
  assign pp_15_34 = ~(be_2x_15_4 & be_x_15_4);
  assign pp_15_35 = ~(be_2x_15_5 & be_x_15_5);
  assign pp_15_36 = ~(be_2x_15_6 & be_x_15_6);
  assign pp_15_37 = ~(be_2x_15_7 & be_x_15_7);
  assign pp_15_38 = ~(be_2x_15_8 & be_x_15_8);
  assign pp_15_39 = ~(be_2x_15_9 & be_x_15_9);
  assign pp_15_40 = ~(be_2x_15_10 & be_x_15_10);
  assign pp_15_41 = ~(be_2x_15_11 & be_x_15_11);
  assign pp_15_42 = ~(be_2x_15_12 & be_x_15_12);
  assign pp_15_43 = ~(be_2x_15_13 & be_x_15_13);
  assign pp_15_44 = ~(be_2x_15_14 & be_x_15_14);
  assign pp_15_45 = ~(be_2x_15_15 & be_x_15_15);
  assign pp_15_46 = ~(be_2x_15_16 & be_x_15_16);
  assign pp_15_47 = ~(be_2x_15_17 & be_x_15_17);
  assign pp_15_48 = ~(be_2x_15_18 & be_x_15_18);
  assign pp_15_49 = ~(be_2x_15_19 & be_x_15_19);
  assign pp_15_50 = ~(be_2x_15_20 & be_x_15_20);
  assign pp_15_51 = ~(be_2x_15_21 & be_x_15_21);
  assign pp_15_52 = ~(be_2x_15_22 & be_x_15_22);
  assign pp_15_53 = ~(be_2x_15_23 & be_x_15_23);
  assign pp_15_54 = ~(be_2x_15_24 & be_x_15_24);
  assign pp_15_55 = ~(be_2x_15_25 & be_x_15_25);
  assign pp_15_56 = ~(be_2x_15_26 & be_x_15_26);
  assign pp_15_57 = ~(be_2x_15_27 & be_x_15_27);
  assign pp_15_58 = ~(be_2x_15_28 & be_x_15_28);
  assign pp_15_59 = ~(be_2x_15_29 & be_x_15_29);
  assign pp_15_60 = ~(be_2x_15_30 & be_x_15_30);
  assign pp_15_61 = ~(be_2x_15_31 & be_x_15_31);
  assign pp_15_62 = ~(be_2x_15_32 & be_x_15_32);
  assign pp_15_63 = ~(be_2x_15_33 & be_x_15_33);
  assign pp_16_32 = ~(be_2x_16_0 & be_x_16_0);
  assign pp_16_33 = ~(be_2x_16_1 & be_x_16_1);
  assign pp_16_34 = ~(be_2x_16_2 & be_x_16_2);
  assign pp_16_35 = ~(be_2x_16_3 & be_x_16_3);
  assign pp_16_36 = ~(be_2x_16_4 & be_x_16_4);
  assign pp_16_37 = ~(be_2x_16_5 & be_x_16_5);
  assign pp_16_38 = ~(be_2x_16_6 & be_x_16_6);
  assign pp_16_39 = ~(be_2x_16_7 & be_x_16_7);
  assign pp_16_40 = ~(be_2x_16_8 & be_x_16_8);
  assign pp_16_41 = ~(be_2x_16_9 & be_x_16_9);
  assign pp_16_42 = ~(be_2x_16_10 & be_x_16_10);
  assign pp_16_43 = ~(be_2x_16_11 & be_x_16_11);
  assign pp_16_44 = ~(be_2x_16_12 & be_x_16_12);
  assign pp_16_45 = ~(be_2x_16_13 & be_x_16_13);
  assign pp_16_46 = ~(be_2x_16_14 & be_x_16_14);
  assign pp_16_47 = ~(be_2x_16_15 & be_x_16_15);
  assign pp_16_48 = ~(be_2x_16_16 & be_x_16_16);
  assign pp_16_49 = ~(be_2x_16_17 & be_x_16_17);
  assign pp_16_50 = ~(be_2x_16_18 & be_x_16_18);
  assign pp_16_51 = ~(be_2x_16_19 & be_x_16_19);
  assign pp_16_52 = ~(be_2x_16_20 & be_x_16_20);
  assign pp_16_53 = ~(be_2x_16_21 & be_x_16_21);
  assign pp_16_54 = ~(be_2x_16_22 & be_x_16_22);
  assign pp_16_55 = ~(be_2x_16_23 & be_x_16_23);
  assign pp_16_56 = ~(be_2x_16_24 & be_x_16_24);
  assign pp_16_57 = ~(be_2x_16_25 & be_x_16_25);
  assign pp_16_58 = ~(be_2x_16_26 & be_x_16_26);
  assign pp_16_59 = ~(be_2x_16_27 & be_x_16_27);
  assign pp_16_60 = ~(be_2x_16_28 & be_x_16_28);
  assign pp_16_61 = ~(be_2x_16_29 & be_x_16_29);
  assign pp_16_62 = ~(be_2x_16_30 & be_x_16_30);
  assign pp_16_63 = ~(be_2x_16_31 & be_x_16_31);
  assign pp_1_10 = ~(be_2x_1_8 & be_x_1_8);
  assign pp_1_11 = ~(be_2x_1_9 & be_x_1_9);
  assign pp_1_12 = ~(be_2x_1_10 & be_x_1_10);
  assign pp_1_13 = ~(be_2x_1_11 & be_x_1_11);
  assign pp_1_14 = ~(be_2x_1_12 & be_x_1_12);
  assign pp_1_15 = ~(be_2x_1_13 & be_x_1_13);
  assign pp_1_16 = ~(be_2x_1_14 & be_x_1_14);
  assign pp_1_17 = ~(be_2x_1_15 & be_x_1_15);
  assign pp_1_18 = ~(be_2x_1_16 & be_x_1_16);
  assign pp_1_19 = ~(be_2x_1_17 & be_x_1_17);
  assign pp_1_2 = ~(be_2x_1_0 & be_x_1_0);
  assign pp_1_20 = ~(be_2x_1_18 & be_x_1_18);
  assign pp_1_21 = ~(be_2x_1_19 & be_x_1_19);
  assign pp_1_22 = ~(be_2x_1_20 & be_x_1_20);
  assign pp_1_23 = ~(be_2x_1_21 & be_x_1_21);
  assign pp_1_24 = ~(be_2x_1_22 & be_x_1_22);
  assign pp_1_25 = ~(be_2x_1_23 & be_x_1_23);
  assign pp_1_26 = ~(be_2x_1_24 & be_x_1_24);
  assign pp_1_27 = ~(be_2x_1_25 & be_x_1_25);
  assign pp_1_28 = ~(be_2x_1_26 & be_x_1_26);
  assign pp_1_29 = ~(be_2x_1_27 & be_x_1_27);
  assign pp_1_3 = ~(be_2x_1_1 & be_x_1_1);
  assign pp_1_30 = ~(be_2x_1_28 & be_x_1_28);
  assign pp_1_31 = ~(be_2x_1_29 & be_x_1_29);
  assign pp_1_32 = ~(be_2x_1_30 & be_x_1_30);
  assign pp_1_33 = ~(be_2x_1_31 & be_x_1_31);
  assign pp_1_34 = ~(be_2x_1_32 & be_x_1_32);
  assign pp_1_35 = ~(be_2x_1_33 & be_x_1_33);
  assign pp_1_4 = ~(be_2x_1_2 & be_x_1_2);
  assign pp_1_5 = ~(be_2x_1_3 & be_x_1_3);
  assign pp_1_6 = ~(be_2x_1_4 & be_x_1_4);
  assign pp_1_7 = ~(be_2x_1_5 & be_x_1_5);
  assign pp_1_8 = ~(be_2x_1_6 & be_x_1_6);
  assign pp_1_9 = ~(be_2x_1_7 & be_x_1_7);
  assign pp_2_10 = ~(be_2x_2_6 & be_x_2_6);
  assign pp_2_11 = ~(be_2x_2_7 & be_x_2_7);
  assign pp_2_12 = ~(be_2x_2_8 & be_x_2_8);
  assign pp_2_13 = ~(be_2x_2_9 & be_x_2_9);
  assign pp_2_14 = ~(be_2x_2_10 & be_x_2_10);
  assign pp_2_15 = ~(be_2x_2_11 & be_x_2_11);
  assign pp_2_16 = ~(be_2x_2_12 & be_x_2_12);
  assign pp_2_17 = ~(be_2x_2_13 & be_x_2_13);
  assign pp_2_18 = ~(be_2x_2_14 & be_x_2_14);
  assign pp_2_19 = ~(be_2x_2_15 & be_x_2_15);
  assign pp_2_20 = ~(be_2x_2_16 & be_x_2_16);
  assign pp_2_21 = ~(be_2x_2_17 & be_x_2_17);
  assign pp_2_22 = ~(be_2x_2_18 & be_x_2_18);
  assign pp_2_23 = ~(be_2x_2_19 & be_x_2_19);
  assign pp_2_24 = ~(be_2x_2_20 & be_x_2_20);
  assign pp_2_25 = ~(be_2x_2_21 & be_x_2_21);
  assign pp_2_26 = ~(be_2x_2_22 & be_x_2_22);
  assign pp_2_27 = ~(be_2x_2_23 & be_x_2_23);
  assign pp_2_28 = ~(be_2x_2_24 & be_x_2_24);
  assign pp_2_29 = ~(be_2x_2_25 & be_x_2_25);
  assign pp_2_30 = ~(be_2x_2_26 & be_x_2_26);
  assign pp_2_31 = ~(be_2x_2_27 & be_x_2_27);
  assign pp_2_32 = ~(be_2x_2_28 & be_x_2_28);
  assign pp_2_33 = ~(be_2x_2_29 & be_x_2_29);
  assign pp_2_34 = ~(be_2x_2_30 & be_x_2_30);
  assign pp_2_35 = ~(be_2x_2_31 & be_x_2_31);
  assign pp_2_36 = ~(be_2x_2_32 & be_x_2_32);
  assign pp_2_37 = ~(be_2x_2_33 & be_x_2_33);
  assign pp_2_4 = ~(be_2x_2_0 & be_x_2_0);
  assign pp_2_5 = ~(be_2x_2_1 & be_x_2_1);
  assign pp_2_6 = ~(be_2x_2_2 & be_x_2_2);
  assign pp_2_7 = ~(be_2x_2_3 & be_x_2_3);
  assign pp_2_8 = ~(be_2x_2_4 & be_x_2_4);
  assign pp_2_9 = ~(be_2x_2_5 & be_x_2_5);
  assign pp_3_10 = ~(be_2x_3_4 & be_x_3_4);
  assign pp_3_11 = ~(be_2x_3_5 & be_x_3_5);
  assign pp_3_12 = ~(be_2x_3_6 & be_x_3_6);
  assign pp_3_13 = ~(be_2x_3_7 & be_x_3_7);
  assign pp_3_14 = ~(be_2x_3_8 & be_x_3_8);
  assign pp_3_15 = ~(be_2x_3_9 & be_x_3_9);
  assign pp_3_16 = ~(be_2x_3_10 & be_x_3_10);
  assign pp_3_17 = ~(be_2x_3_11 & be_x_3_11);
  assign pp_3_18 = ~(be_2x_3_12 & be_x_3_12);
  assign pp_3_19 = ~(be_2x_3_13 & be_x_3_13);
  assign pp_3_20 = ~(be_2x_3_14 & be_x_3_14);
  assign pp_3_21 = ~(be_2x_3_15 & be_x_3_15);
  assign pp_3_22 = ~(be_2x_3_16 & be_x_3_16);
  assign pp_3_23 = ~(be_2x_3_17 & be_x_3_17);
  assign pp_3_24 = ~(be_2x_3_18 & be_x_3_18);
  assign pp_3_25 = ~(be_2x_3_19 & be_x_3_19);
  assign pp_3_26 = ~(be_2x_3_20 & be_x_3_20);
  assign pp_3_27 = ~(be_2x_3_21 & be_x_3_21);
  assign pp_3_28 = ~(be_2x_3_22 & be_x_3_22);
  assign pp_3_29 = ~(be_2x_3_23 & be_x_3_23);
  assign pp_3_30 = ~(be_2x_3_24 & be_x_3_24);
  assign pp_3_31 = ~(be_2x_3_25 & be_x_3_25);
  assign pp_3_32 = ~(be_2x_3_26 & be_x_3_26);
  assign pp_3_33 = ~(be_2x_3_27 & be_x_3_27);
  assign pp_3_34 = ~(be_2x_3_28 & be_x_3_28);
  assign pp_3_35 = ~(be_2x_3_29 & be_x_3_29);
  assign pp_3_36 = ~(be_2x_3_30 & be_x_3_30);
  assign pp_3_37 = ~(be_2x_3_31 & be_x_3_31);
  assign pp_3_38 = ~(be_2x_3_32 & be_x_3_32);
  assign pp_3_39 = ~(be_2x_3_33 & be_x_3_33);
  assign pp_3_6 = ~(be_2x_3_0 & be_x_3_0);
  assign pp_3_7 = ~(be_2x_3_1 & be_x_3_1);
  assign pp_3_8 = ~(be_2x_3_2 & be_x_3_2);
  assign pp_3_9 = ~(be_2x_3_3 & be_x_3_3);
  assign pp_4_10 = ~(be_2x_4_2 & be_x_4_2);
  assign pp_4_11 = ~(be_2x_4_3 & be_x_4_3);
  assign pp_4_12 = ~(be_2x_4_4 & be_x_4_4);
  assign pp_4_13 = ~(be_2x_4_5 & be_x_4_5);
  assign pp_4_14 = ~(be_2x_4_6 & be_x_4_6);
  assign pp_4_15 = ~(be_2x_4_7 & be_x_4_7);
  assign pp_4_16 = ~(be_2x_4_8 & be_x_4_8);
  assign pp_4_17 = ~(be_2x_4_9 & be_x_4_9);
  assign pp_4_18 = ~(be_2x_4_10 & be_x_4_10);
  assign pp_4_19 = ~(be_2x_4_11 & be_x_4_11);
  assign pp_4_20 = ~(be_2x_4_12 & be_x_4_12);
  assign pp_4_21 = ~(be_2x_4_13 & be_x_4_13);
  assign pp_4_22 = ~(be_2x_4_14 & be_x_4_14);
  assign pp_4_23 = ~(be_2x_4_15 & be_x_4_15);
  assign pp_4_24 = ~(be_2x_4_16 & be_x_4_16);
  assign pp_4_25 = ~(be_2x_4_17 & be_x_4_17);
  assign pp_4_26 = ~(be_2x_4_18 & be_x_4_18);
  assign pp_4_27 = ~(be_2x_4_19 & be_x_4_19);
  assign pp_4_28 = ~(be_2x_4_20 & be_x_4_20);
  assign pp_4_29 = ~(be_2x_4_21 & be_x_4_21);
  assign pp_4_30 = ~(be_2x_4_22 & be_x_4_22);
  assign pp_4_31 = ~(be_2x_4_23 & be_x_4_23);
  assign pp_4_32 = ~(be_2x_4_24 & be_x_4_24);
  assign pp_4_33 = ~(be_2x_4_25 & be_x_4_25);
  assign pp_4_34 = ~(be_2x_4_26 & be_x_4_26);
  assign pp_4_35 = ~(be_2x_4_27 & be_x_4_27);
  assign pp_4_36 = ~(be_2x_4_28 & be_x_4_28);
  assign pp_4_37 = ~(be_2x_4_29 & be_x_4_29);
  assign pp_4_38 = ~(be_2x_4_30 & be_x_4_30);
  assign pp_4_39 = ~(be_2x_4_31 & be_x_4_31);
  assign pp_4_40 = ~(be_2x_4_32 & be_x_4_32);
  assign pp_4_41 = ~(be_2x_4_33 & be_x_4_33);
  assign pp_4_8 = ~(be_2x_4_0 & be_x_4_0);
  assign pp_4_9 = ~(be_2x_4_1 & be_x_4_1);
  assign pp_5_10 = ~(be_2x_5_0 & be_x_5_0);
  assign pp_5_11 = ~(be_2x_5_1 & be_x_5_1);
  assign pp_5_12 = ~(be_2x_5_2 & be_x_5_2);
  assign pp_5_13 = ~(be_2x_5_3 & be_x_5_3);
  assign pp_5_14 = ~(be_2x_5_4 & be_x_5_4);
  assign pp_5_15 = ~(be_2x_5_5 & be_x_5_5);
  assign pp_5_16 = ~(be_2x_5_6 & be_x_5_6);
  assign pp_5_17 = ~(be_2x_5_7 & be_x_5_7);
  assign pp_5_18 = ~(be_2x_5_8 & be_x_5_8);
  assign pp_5_19 = ~(be_2x_5_9 & be_x_5_9);
  assign pp_5_20 = ~(be_2x_5_10 & be_x_5_10);
  assign pp_5_21 = ~(be_2x_5_11 & be_x_5_11);
  assign pp_5_22 = ~(be_2x_5_12 & be_x_5_12);
  assign pp_5_23 = ~(be_2x_5_13 & be_x_5_13);
  assign pp_5_24 = ~(be_2x_5_14 & be_x_5_14);
  assign pp_5_25 = ~(be_2x_5_15 & be_x_5_15);
  assign pp_5_26 = ~(be_2x_5_16 & be_x_5_16);
  assign pp_5_27 = ~(be_2x_5_17 & be_x_5_17);
  assign pp_5_28 = ~(be_2x_5_18 & be_x_5_18);
  assign pp_5_29 = ~(be_2x_5_19 & be_x_5_19);
  assign pp_5_30 = ~(be_2x_5_20 & be_x_5_20);
  assign pp_5_31 = ~(be_2x_5_21 & be_x_5_21);
  assign pp_5_32 = ~(be_2x_5_22 & be_x_5_22);
  assign pp_5_33 = ~(be_2x_5_23 & be_x_5_23);
  assign pp_5_34 = ~(be_2x_5_24 & be_x_5_24);
  assign pp_5_35 = ~(be_2x_5_25 & be_x_5_25);
  assign pp_5_36 = ~(be_2x_5_26 & be_x_5_26);
  assign pp_5_37 = ~(be_2x_5_27 & be_x_5_27);
  assign pp_5_38 = ~(be_2x_5_28 & be_x_5_28);
  assign pp_5_39 = ~(be_2x_5_29 & be_x_5_29);
  assign pp_5_40 = ~(be_2x_5_30 & be_x_5_30);
  assign pp_5_41 = ~(be_2x_5_31 & be_x_5_31);
  assign pp_5_42 = ~(be_2x_5_32 & be_x_5_32);
  assign pp_5_43 = ~(be_2x_5_33 & be_x_5_33);
  assign pp_6_12 = ~(be_2x_6_0 & be_x_6_0);
  assign pp_6_13 = ~(be_2x_6_1 & be_x_6_1);
  assign pp_6_14 = ~(be_2x_6_2 & be_x_6_2);
  assign pp_6_15 = ~(be_2x_6_3 & be_x_6_3);
  assign pp_6_16 = ~(be_2x_6_4 & be_x_6_4);
  assign pp_6_17 = ~(be_2x_6_5 & be_x_6_5);
  assign pp_6_18 = ~(be_2x_6_6 & be_x_6_6);
  assign pp_6_19 = ~(be_2x_6_7 & be_x_6_7);
  assign pp_6_20 = ~(be_2x_6_8 & be_x_6_8);
  assign pp_6_21 = ~(be_2x_6_9 & be_x_6_9);
  assign pp_6_22 = ~(be_2x_6_10 & be_x_6_10);
  assign pp_6_23 = ~(be_2x_6_11 & be_x_6_11);
  assign pp_6_24 = ~(be_2x_6_12 & be_x_6_12);
  assign pp_6_25 = ~(be_2x_6_13 & be_x_6_13);
  assign pp_6_26 = ~(be_2x_6_14 & be_x_6_14);
  assign pp_6_27 = ~(be_2x_6_15 & be_x_6_15);
  assign pp_6_28 = ~(be_2x_6_16 & be_x_6_16);
  assign pp_6_29 = ~(be_2x_6_17 & be_x_6_17);
  assign pp_6_30 = ~(be_2x_6_18 & be_x_6_18);
  assign pp_6_31 = ~(be_2x_6_19 & be_x_6_19);
  assign pp_6_32 = ~(be_2x_6_20 & be_x_6_20);
  assign pp_6_33 = ~(be_2x_6_21 & be_x_6_21);
  assign pp_6_34 = ~(be_2x_6_22 & be_x_6_22);
  assign pp_6_35 = ~(be_2x_6_23 & be_x_6_23);
  assign pp_6_36 = ~(be_2x_6_24 & be_x_6_24);
  assign pp_6_37 = ~(be_2x_6_25 & be_x_6_25);
  assign pp_6_38 = ~(be_2x_6_26 & be_x_6_26);
  assign pp_6_39 = ~(be_2x_6_27 & be_x_6_27);
  assign pp_6_40 = ~(be_2x_6_28 & be_x_6_28);
  assign pp_6_41 = ~(be_2x_6_29 & be_x_6_29);
  assign pp_6_42 = ~(be_2x_6_30 & be_x_6_30);
  assign pp_6_43 = ~(be_2x_6_31 & be_x_6_31);
  assign pp_6_44 = ~(be_2x_6_32 & be_x_6_32);
  assign pp_6_45 = ~(be_2x_6_33 & be_x_6_33);
  assign pp_7_14 = ~(be_2x_7_0 & be_x_7_0);
  assign pp_7_15 = ~(be_2x_7_1 & be_x_7_1);
  assign pp_7_16 = ~(be_2x_7_2 & be_x_7_2);
  assign pp_7_17 = ~(be_2x_7_3 & be_x_7_3);
  assign pp_7_18 = ~(be_2x_7_4 & be_x_7_4);
  assign pp_7_19 = ~(be_2x_7_5 & be_x_7_5);
  assign pp_7_20 = ~(be_2x_7_6 & be_x_7_6);
  assign pp_7_21 = ~(be_2x_7_7 & be_x_7_7);
  assign pp_7_22 = ~(be_2x_7_8 & be_x_7_8);
  assign pp_7_23 = ~(be_2x_7_9 & be_x_7_9);
  assign pp_7_24 = ~(be_2x_7_10 & be_x_7_10);
  assign pp_7_25 = ~(be_2x_7_11 & be_x_7_11);
  assign pp_7_26 = ~(be_2x_7_12 & be_x_7_12);
  assign pp_7_27 = ~(be_2x_7_13 & be_x_7_13);
  assign pp_7_28 = ~(be_2x_7_14 & be_x_7_14);
  assign pp_7_29 = ~(be_2x_7_15 & be_x_7_15);
  assign pp_7_30 = ~(be_2x_7_16 & be_x_7_16);
  assign pp_7_31 = ~(be_2x_7_17 & be_x_7_17);
  assign pp_7_32 = ~(be_2x_7_18 & be_x_7_18);
  assign pp_7_33 = ~(be_2x_7_19 & be_x_7_19);
  assign pp_7_34 = ~(be_2x_7_20 & be_x_7_20);
  assign pp_7_35 = ~(be_2x_7_21 & be_x_7_21);
  assign pp_7_36 = ~(be_2x_7_22 & be_x_7_22);
  assign pp_7_37 = ~(be_2x_7_23 & be_x_7_23);
  assign pp_7_38 = ~(be_2x_7_24 & be_x_7_24);
  assign pp_7_39 = ~(be_2x_7_25 & be_x_7_25);
  assign pp_7_40 = ~(be_2x_7_26 & be_x_7_26);
  assign pp_7_41 = ~(be_2x_7_27 & be_x_7_27);
  assign pp_7_42 = ~(be_2x_7_28 & be_x_7_28);
  assign pp_7_43 = ~(be_2x_7_29 & be_x_7_29);
  assign pp_7_44 = ~(be_2x_7_30 & be_x_7_30);
  assign pp_7_45 = ~(be_2x_7_31 & be_x_7_31);
  assign pp_7_46 = ~(be_2x_7_32 & be_x_7_32);
  assign pp_7_47 = ~(be_2x_7_33 & be_x_7_33);
  assign pp_8_16 = ~(be_2x_8_0 & be_x_8_0);
  assign pp_8_17 = ~(be_2x_8_1 & be_x_8_1);
  assign pp_8_18 = ~(be_2x_8_2 & be_x_8_2);
  assign pp_8_19 = ~(be_2x_8_3 & be_x_8_3);
  assign pp_8_20 = ~(be_2x_8_4 & be_x_8_4);
  assign pp_8_21 = ~(be_2x_8_5 & be_x_8_5);
  assign pp_8_22 = ~(be_2x_8_6 & be_x_8_6);
  assign pp_8_23 = ~(be_2x_8_7 & be_x_8_7);
  assign pp_8_24 = ~(be_2x_8_8 & be_x_8_8);
  assign pp_8_25 = ~(be_2x_8_9 & be_x_8_9);
  assign pp_8_26 = ~(be_2x_8_10 & be_x_8_10);
  assign pp_8_27 = ~(be_2x_8_11 & be_x_8_11);
  assign pp_8_28 = ~(be_2x_8_12 & be_x_8_12);
  assign pp_8_29 = ~(be_2x_8_13 & be_x_8_13);
  assign pp_8_30 = ~(be_2x_8_14 & be_x_8_14);
  assign pp_8_31 = ~(be_2x_8_15 & be_x_8_15);
  assign pp_8_32 = ~(be_2x_8_16 & be_x_8_16);
  assign pp_8_33 = ~(be_2x_8_17 & be_x_8_17);
  assign pp_8_34 = ~(be_2x_8_18 & be_x_8_18);
  assign pp_8_35 = ~(be_2x_8_19 & be_x_8_19);
  assign pp_8_36 = ~(be_2x_8_20 & be_x_8_20);
  assign pp_8_37 = ~(be_2x_8_21 & be_x_8_21);
  assign pp_8_38 = ~(be_2x_8_22 & be_x_8_22);
  assign pp_8_39 = ~(be_2x_8_23 & be_x_8_23);
  assign pp_8_40 = ~(be_2x_8_24 & be_x_8_24);
  assign pp_8_41 = ~(be_2x_8_25 & be_x_8_25);
  assign pp_8_42 = ~(be_2x_8_26 & be_x_8_26);
  assign pp_8_43 = ~(be_2x_8_27 & be_x_8_27);
  assign pp_8_44 = ~(be_2x_8_28 & be_x_8_28);
  assign pp_8_45 = ~(be_2x_8_29 & be_x_8_29);
  assign pp_8_46 = ~(be_2x_8_30 & be_x_8_30);
  assign pp_8_47 = ~(be_2x_8_31 & be_x_8_31);
  assign pp_8_48 = ~(be_2x_8_32 & be_x_8_32);
  assign pp_8_49 = ~(be_2x_8_33 & be_x_8_33);
  assign pp_9_18 = ~(be_2x_9_0 & be_x_9_0);
  assign pp_9_19 = ~(be_2x_9_1 & be_x_9_1);
  assign pp_9_20 = ~(be_2x_9_2 & be_x_9_2);
  assign pp_9_21 = ~(be_2x_9_3 & be_x_9_3);
  assign pp_9_22 = ~(be_2x_9_4 & be_x_9_4);
  assign pp_9_23 = ~(be_2x_9_5 & be_x_9_5);
  assign pp_9_24 = ~(be_2x_9_6 & be_x_9_6);
  assign pp_9_25 = ~(be_2x_9_7 & be_x_9_7);
  assign pp_9_26 = ~(be_2x_9_8 & be_x_9_8);
  assign pp_9_27 = ~(be_2x_9_9 & be_x_9_9);
  assign pp_9_28 = ~(be_2x_9_10 & be_x_9_10);
  assign pp_9_29 = ~(be_2x_9_11 & be_x_9_11);
  assign pp_9_30 = ~(be_2x_9_12 & be_x_9_12);
  assign pp_9_31 = ~(be_2x_9_13 & be_x_9_13);
  assign pp_9_32 = ~(be_2x_9_14 & be_x_9_14);
  assign pp_9_33 = ~(be_2x_9_15 & be_x_9_15);
  assign pp_9_34 = ~(be_2x_9_16 & be_x_9_16);
  assign pp_9_35 = ~(be_2x_9_17 & be_x_9_17);
  assign pp_9_36 = ~(be_2x_9_18 & be_x_9_18);
  assign pp_9_37 = ~(be_2x_9_19 & be_x_9_19);
  assign pp_9_38 = ~(be_2x_9_20 & be_x_9_20);
  assign pp_9_39 = ~(be_2x_9_21 & be_x_9_21);
  assign pp_9_40 = ~(be_2x_9_22 & be_x_9_22);
  assign pp_9_41 = ~(be_2x_9_23 & be_x_9_23);
  assign pp_9_42 = ~(be_2x_9_24 & be_x_9_24);
  assign pp_9_43 = ~(be_2x_9_25 & be_x_9_25);
  assign pp_9_44 = ~(be_2x_9_26 & be_x_9_26);
  assign pp_9_45 = ~(be_2x_9_27 & be_x_9_27);
  assign pp_9_46 = ~(be_2x_9_28 & be_x_9_28);
  assign pp_9_47 = ~(be_2x_9_29 & be_x_9_29);
  assign pp_9_48 = ~(be_2x_9_30 & be_x_9_30);
  assign pp_9_49 = ~(be_2x_9_31 & be_x_9_31);
  assign pp_9_50 = ~(be_2x_9_32 & be_x_9_32);
  assign pp_9_51 = ~(be_2x_9_33 & be_x_9_33);
  assign px_0_0 = be_neg_0;
  assign px_0_1 = be_neg_0 ^ x_0;
  assign px_0_10 = be_neg_0 ^ x_9;
  assign px_0_11 = be_neg_0 ^ x_10;
  assign px_0_12 = be_neg_0 ^ x_11;
  assign px_0_13 = be_neg_0 ^ x_12;
  assign px_0_14 = be_neg_0 ^ x_13;
  assign px_0_15 = be_neg_0 ^ x_14;
  assign px_0_16 = be_neg_0 ^ x_15;
  assign px_0_17 = be_neg_0 ^ x_16;
  assign px_0_18 = be_neg_0 ^ x_17;
  assign px_0_19 = be_neg_0 ^ x_18;
  assign px_0_2 = be_neg_0 ^ x_1;
  assign px_0_20 = be_neg_0 ^ x_19;
  assign px_0_21 = be_neg_0 ^ x_20;
  assign px_0_22 = be_neg_0 ^ x_21;
  assign px_0_23 = be_neg_0 ^ x_22;
  assign px_0_24 = be_neg_0 ^ x_23;
  assign px_0_25 = be_neg_0 ^ x_24;
  assign px_0_26 = be_neg_0 ^ x_25;
  assign px_0_27 = be_neg_0 ^ x_26;
  assign px_0_28 = be_neg_0 ^ x_27;
  assign px_0_29 = be_neg_0 ^ x_28;
  assign px_0_3 = be_neg_0 ^ x_2;
  assign px_0_30 = be_neg_0 ^ x_29;
  assign px_0_31 = be_neg_0 ^ x_30;
  assign px_0_32 = be_neg_0 ^ x_31;
  assign px_0_33 = be_neg_0 ^ zero;
  assign px_0_34 = be_neg_0 ^ zero;
  assign px_0_4 = be_neg_0 ^ x_3;
  assign px_0_5 = be_neg_0 ^ x_4;
  assign px_0_6 = be_neg_0 ^ x_5;
  assign px_0_7 = be_neg_0 ^ x_6;
  assign px_0_8 = be_neg_0 ^ x_7;
  assign px_0_9 = be_neg_0 ^ x_8;
  assign px_10_0 = be_neg_10;
  assign px_10_1 = be_neg_10 ^ x_0;
  assign px_10_10 = be_neg_10 ^ x_9;
  assign px_10_11 = be_neg_10 ^ x_10;
  assign px_10_12 = be_neg_10 ^ x_11;
  assign px_10_13 = be_neg_10 ^ x_12;
  assign px_10_14 = be_neg_10 ^ x_13;
  assign px_10_15 = be_neg_10 ^ x_14;
  assign px_10_16 = be_neg_10 ^ x_15;
  assign px_10_17 = be_neg_10 ^ x_16;
  assign px_10_18 = be_neg_10 ^ x_17;
  assign px_10_19 = be_neg_10 ^ x_18;
  assign px_10_2 = be_neg_10 ^ x_1;
  assign px_10_20 = be_neg_10 ^ x_19;
  assign px_10_21 = be_neg_10 ^ x_20;
  assign px_10_22 = be_neg_10 ^ x_21;
  assign px_10_23 = be_neg_10 ^ x_22;
  assign px_10_24 = be_neg_10 ^ x_23;
  assign px_10_25 = be_neg_10 ^ x_24;
  assign px_10_26 = be_neg_10 ^ x_25;
  assign px_10_27 = be_neg_10 ^ x_26;
  assign px_10_28 = be_neg_10 ^ x_27;
  assign px_10_29 = be_neg_10 ^ x_28;
  assign px_10_3 = be_neg_10 ^ x_2;
  assign px_10_30 = be_neg_10 ^ x_29;
  assign px_10_31 = be_neg_10 ^ x_30;
  assign px_10_32 = be_neg_10 ^ x_31;
  assign px_10_33 = be_neg_10 ^ zero;
  assign px_10_34 = be_neg_10 ^ zero;
  assign px_10_4 = be_neg_10 ^ x_3;
  assign px_10_5 = be_neg_10 ^ x_4;
  assign px_10_6 = be_neg_10 ^ x_5;
  assign px_10_7 = be_neg_10 ^ x_6;
  assign px_10_8 = be_neg_10 ^ x_7;
  assign px_10_9 = be_neg_10 ^ x_8;
  assign px_11_0 = be_neg_11;
  assign px_11_1 = be_neg_11 ^ x_0;
  assign px_11_10 = be_neg_11 ^ x_9;
  assign px_11_11 = be_neg_11 ^ x_10;
  assign px_11_12 = be_neg_11 ^ x_11;
  assign px_11_13 = be_neg_11 ^ x_12;
  assign px_11_14 = be_neg_11 ^ x_13;
  assign px_11_15 = be_neg_11 ^ x_14;
  assign px_11_16 = be_neg_11 ^ x_15;
  assign px_11_17 = be_neg_11 ^ x_16;
  assign px_11_18 = be_neg_11 ^ x_17;
  assign px_11_19 = be_neg_11 ^ x_18;
  assign px_11_2 = be_neg_11 ^ x_1;
  assign px_11_20 = be_neg_11 ^ x_19;
  assign px_11_21 = be_neg_11 ^ x_20;
  assign px_11_22 = be_neg_11 ^ x_21;
  assign px_11_23 = be_neg_11 ^ x_22;
  assign px_11_24 = be_neg_11 ^ x_23;
  assign px_11_25 = be_neg_11 ^ x_24;
  assign px_11_26 = be_neg_11 ^ x_25;
  assign px_11_27 = be_neg_11 ^ x_26;
  assign px_11_28 = be_neg_11 ^ x_27;
  assign px_11_29 = be_neg_11 ^ x_28;
  assign px_11_3 = be_neg_11 ^ x_2;
  assign px_11_30 = be_neg_11 ^ x_29;
  assign px_11_31 = be_neg_11 ^ x_30;
  assign px_11_32 = be_neg_11 ^ x_31;
  assign px_11_33 = be_neg_11 ^ zero;
  assign px_11_34 = be_neg_11 ^ zero;
  assign px_11_4 = be_neg_11 ^ x_3;
  assign px_11_5 = be_neg_11 ^ x_4;
  assign px_11_6 = be_neg_11 ^ x_5;
  assign px_11_7 = be_neg_11 ^ x_6;
  assign px_11_8 = be_neg_11 ^ x_7;
  assign px_11_9 = be_neg_11 ^ x_8;
  assign px_12_0 = be_neg_12;
  assign px_12_1 = be_neg_12 ^ x_0;
  assign px_12_10 = be_neg_12 ^ x_9;
  assign px_12_11 = be_neg_12 ^ x_10;
  assign px_12_12 = be_neg_12 ^ x_11;
  assign px_12_13 = be_neg_12 ^ x_12;
  assign px_12_14 = be_neg_12 ^ x_13;
  assign px_12_15 = be_neg_12 ^ x_14;
  assign px_12_16 = be_neg_12 ^ x_15;
  assign px_12_17 = be_neg_12 ^ x_16;
  assign px_12_18 = be_neg_12 ^ x_17;
  assign px_12_19 = be_neg_12 ^ x_18;
  assign px_12_2 = be_neg_12 ^ x_1;
  assign px_12_20 = be_neg_12 ^ x_19;
  assign px_12_21 = be_neg_12 ^ x_20;
  assign px_12_22 = be_neg_12 ^ x_21;
  assign px_12_23 = be_neg_12 ^ x_22;
  assign px_12_24 = be_neg_12 ^ x_23;
  assign px_12_25 = be_neg_12 ^ x_24;
  assign px_12_26 = be_neg_12 ^ x_25;
  assign px_12_27 = be_neg_12 ^ x_26;
  assign px_12_28 = be_neg_12 ^ x_27;
  assign px_12_29 = be_neg_12 ^ x_28;
  assign px_12_3 = be_neg_12 ^ x_2;
  assign px_12_30 = be_neg_12 ^ x_29;
  assign px_12_31 = be_neg_12 ^ x_30;
  assign px_12_32 = be_neg_12 ^ x_31;
  assign px_12_33 = be_neg_12 ^ zero;
  assign px_12_34 = be_neg_12 ^ zero;
  assign px_12_4 = be_neg_12 ^ x_3;
  assign px_12_5 = be_neg_12 ^ x_4;
  assign px_12_6 = be_neg_12 ^ x_5;
  assign px_12_7 = be_neg_12 ^ x_6;
  assign px_12_8 = be_neg_12 ^ x_7;
  assign px_12_9 = be_neg_12 ^ x_8;
  assign px_13_0 = be_neg_13;
  assign px_13_1 = be_neg_13 ^ x_0;
  assign px_13_10 = be_neg_13 ^ x_9;
  assign px_13_11 = be_neg_13 ^ x_10;
  assign px_13_12 = be_neg_13 ^ x_11;
  assign px_13_13 = be_neg_13 ^ x_12;
  assign px_13_14 = be_neg_13 ^ x_13;
  assign px_13_15 = be_neg_13 ^ x_14;
  assign px_13_16 = be_neg_13 ^ x_15;
  assign px_13_17 = be_neg_13 ^ x_16;
  assign px_13_18 = be_neg_13 ^ x_17;
  assign px_13_19 = be_neg_13 ^ x_18;
  assign px_13_2 = be_neg_13 ^ x_1;
  assign px_13_20 = be_neg_13 ^ x_19;
  assign px_13_21 = be_neg_13 ^ x_20;
  assign px_13_22 = be_neg_13 ^ x_21;
  assign px_13_23 = be_neg_13 ^ x_22;
  assign px_13_24 = be_neg_13 ^ x_23;
  assign px_13_25 = be_neg_13 ^ x_24;
  assign px_13_26 = be_neg_13 ^ x_25;
  assign px_13_27 = be_neg_13 ^ x_26;
  assign px_13_28 = be_neg_13 ^ x_27;
  assign px_13_29 = be_neg_13 ^ x_28;
  assign px_13_3 = be_neg_13 ^ x_2;
  assign px_13_30 = be_neg_13 ^ x_29;
  assign px_13_31 = be_neg_13 ^ x_30;
  assign px_13_32 = be_neg_13 ^ x_31;
  assign px_13_33 = be_neg_13 ^ zero;
  assign px_13_34 = be_neg_13 ^ zero;
  assign px_13_4 = be_neg_13 ^ x_3;
  assign px_13_5 = be_neg_13 ^ x_4;
  assign px_13_6 = be_neg_13 ^ x_5;
  assign px_13_7 = be_neg_13 ^ x_6;
  assign px_13_8 = be_neg_13 ^ x_7;
  assign px_13_9 = be_neg_13 ^ x_8;
  assign px_14_0 = be_neg_14;
  assign px_14_1 = be_neg_14 ^ x_0;
  assign px_14_10 = be_neg_14 ^ x_9;
  assign px_14_11 = be_neg_14 ^ x_10;
  assign px_14_12 = be_neg_14 ^ x_11;
  assign px_14_13 = be_neg_14 ^ x_12;
  assign px_14_14 = be_neg_14 ^ x_13;
  assign px_14_15 = be_neg_14 ^ x_14;
  assign px_14_16 = be_neg_14 ^ x_15;
  assign px_14_17 = be_neg_14 ^ x_16;
  assign px_14_18 = be_neg_14 ^ x_17;
  assign px_14_19 = be_neg_14 ^ x_18;
  assign px_14_2 = be_neg_14 ^ x_1;
  assign px_14_20 = be_neg_14 ^ x_19;
  assign px_14_21 = be_neg_14 ^ x_20;
  assign px_14_22 = be_neg_14 ^ x_21;
  assign px_14_23 = be_neg_14 ^ x_22;
  assign px_14_24 = be_neg_14 ^ x_23;
  assign px_14_25 = be_neg_14 ^ x_24;
  assign px_14_26 = be_neg_14 ^ x_25;
  assign px_14_27 = be_neg_14 ^ x_26;
  assign px_14_28 = be_neg_14 ^ x_27;
  assign px_14_29 = be_neg_14 ^ x_28;
  assign px_14_3 = be_neg_14 ^ x_2;
  assign px_14_30 = be_neg_14 ^ x_29;
  assign px_14_31 = be_neg_14 ^ x_30;
  assign px_14_32 = be_neg_14 ^ x_31;
  assign px_14_33 = be_neg_14 ^ zero;
  assign px_14_34 = be_neg_14 ^ zero;
  assign px_14_4 = be_neg_14 ^ x_3;
  assign px_14_5 = be_neg_14 ^ x_4;
  assign px_14_6 = be_neg_14 ^ x_5;
  assign px_14_7 = be_neg_14 ^ x_6;
  assign px_14_8 = be_neg_14 ^ x_7;
  assign px_14_9 = be_neg_14 ^ x_8;
  assign px_15_0 = be_neg_15;
  assign px_15_1 = be_neg_15 ^ x_0;
  assign px_15_10 = be_neg_15 ^ x_9;
  assign px_15_11 = be_neg_15 ^ x_10;
  assign px_15_12 = be_neg_15 ^ x_11;
  assign px_15_13 = be_neg_15 ^ x_12;
  assign px_15_14 = be_neg_15 ^ x_13;
  assign px_15_15 = be_neg_15 ^ x_14;
  assign px_15_16 = be_neg_15 ^ x_15;
  assign px_15_17 = be_neg_15 ^ x_16;
  assign px_15_18 = be_neg_15 ^ x_17;
  assign px_15_19 = be_neg_15 ^ x_18;
  assign px_15_2 = be_neg_15 ^ x_1;
  assign px_15_20 = be_neg_15 ^ x_19;
  assign px_15_21 = be_neg_15 ^ x_20;
  assign px_15_22 = be_neg_15 ^ x_21;
  assign px_15_23 = be_neg_15 ^ x_22;
  assign px_15_24 = be_neg_15 ^ x_23;
  assign px_15_25 = be_neg_15 ^ x_24;
  assign px_15_26 = be_neg_15 ^ x_25;
  assign px_15_27 = be_neg_15 ^ x_26;
  assign px_15_28 = be_neg_15 ^ x_27;
  assign px_15_29 = be_neg_15 ^ x_28;
  assign px_15_3 = be_neg_15 ^ x_2;
  assign px_15_30 = be_neg_15 ^ x_29;
  assign px_15_31 = be_neg_15 ^ x_30;
  assign px_15_32 = be_neg_15 ^ x_31;
  assign px_15_33 = be_neg_15 ^ zero;
  assign px_15_34 = be_neg_15 ^ zero;
  assign px_15_4 = be_neg_15 ^ x_3;
  assign px_15_5 = be_neg_15 ^ x_4;
  assign px_15_6 = be_neg_15 ^ x_5;
  assign px_15_7 = be_neg_15 ^ x_6;
  assign px_15_8 = be_neg_15 ^ x_7;
  assign px_15_9 = be_neg_15 ^ x_8;
  assign px_16_0 = be_neg_16;
  assign px_16_1 = be_neg_16 ^ x_0;
  assign px_16_10 = be_neg_16 ^ x_9;
  assign px_16_11 = be_neg_16 ^ x_10;
  assign px_16_12 = be_neg_16 ^ x_11;
  assign px_16_13 = be_neg_16 ^ x_12;
  assign px_16_14 = be_neg_16 ^ x_13;
  assign px_16_15 = be_neg_16 ^ x_14;
  assign px_16_16 = be_neg_16 ^ x_15;
  assign px_16_17 = be_neg_16 ^ x_16;
  assign px_16_18 = be_neg_16 ^ x_17;
  assign px_16_19 = be_neg_16 ^ x_18;
  assign px_16_2 = be_neg_16 ^ x_1;
  assign px_16_20 = be_neg_16 ^ x_19;
  assign px_16_21 = be_neg_16 ^ x_20;
  assign px_16_22 = be_neg_16 ^ x_21;
  assign px_16_23 = be_neg_16 ^ x_22;
  assign px_16_24 = be_neg_16 ^ x_23;
  assign px_16_25 = be_neg_16 ^ x_24;
  assign px_16_26 = be_neg_16 ^ x_25;
  assign px_16_27 = be_neg_16 ^ x_26;
  assign px_16_28 = be_neg_16 ^ x_27;
  assign px_16_29 = be_neg_16 ^ x_28;
  assign px_16_3 = be_neg_16 ^ x_2;
  assign px_16_30 = be_neg_16 ^ x_29;
  assign px_16_31 = be_neg_16 ^ x_30;
  assign px_16_32 = be_neg_16 ^ x_31;
  assign px_16_33 = be_neg_16 ^ zero;
  assign px_16_34 = be_neg_16 ^ zero;
  assign px_16_4 = be_neg_16 ^ x_3;
  assign px_16_5 = be_neg_16 ^ x_4;
  assign px_16_6 = be_neg_16 ^ x_5;
  assign px_16_7 = be_neg_16 ^ x_6;
  assign px_16_8 = be_neg_16 ^ x_7;
  assign px_16_9 = be_neg_16 ^ x_8;
  assign px_1_0 = be_neg_1;
  assign px_1_1 = be_neg_1 ^ x_0;
  assign px_1_10 = be_neg_1 ^ x_9;
  assign px_1_11 = be_neg_1 ^ x_10;
  assign px_1_12 = be_neg_1 ^ x_11;
  assign px_1_13 = be_neg_1 ^ x_12;
  assign px_1_14 = be_neg_1 ^ x_13;
  assign px_1_15 = be_neg_1 ^ x_14;
  assign px_1_16 = be_neg_1 ^ x_15;
  assign px_1_17 = be_neg_1 ^ x_16;
  assign px_1_18 = be_neg_1 ^ x_17;
  assign px_1_19 = be_neg_1 ^ x_18;
  assign px_1_2 = be_neg_1 ^ x_1;
  assign px_1_20 = be_neg_1 ^ x_19;
  assign px_1_21 = be_neg_1 ^ x_20;
  assign px_1_22 = be_neg_1 ^ x_21;
  assign px_1_23 = be_neg_1 ^ x_22;
  assign px_1_24 = be_neg_1 ^ x_23;
  assign px_1_25 = be_neg_1 ^ x_24;
  assign px_1_26 = be_neg_1 ^ x_25;
  assign px_1_27 = be_neg_1 ^ x_26;
  assign px_1_28 = be_neg_1 ^ x_27;
  assign px_1_29 = be_neg_1 ^ x_28;
  assign px_1_3 = be_neg_1 ^ x_2;
  assign px_1_30 = be_neg_1 ^ x_29;
  assign px_1_31 = be_neg_1 ^ x_30;
  assign px_1_32 = be_neg_1 ^ x_31;
  assign px_1_33 = be_neg_1 ^ zero;
  assign px_1_34 = be_neg_1 ^ zero;
  assign px_1_4 = be_neg_1 ^ x_3;
  assign px_1_5 = be_neg_1 ^ x_4;
  assign px_1_6 = be_neg_1 ^ x_5;
  assign px_1_7 = be_neg_1 ^ x_6;
  assign px_1_8 = be_neg_1 ^ x_7;
  assign px_1_9 = be_neg_1 ^ x_8;
  assign px_2_0 = be_neg_2;
  assign px_2_1 = be_neg_2 ^ x_0;
  assign px_2_10 = be_neg_2 ^ x_9;
  assign px_2_11 = be_neg_2 ^ x_10;
  assign px_2_12 = be_neg_2 ^ x_11;
  assign px_2_13 = be_neg_2 ^ x_12;
  assign px_2_14 = be_neg_2 ^ x_13;
  assign px_2_15 = be_neg_2 ^ x_14;
  assign px_2_16 = be_neg_2 ^ x_15;
  assign px_2_17 = be_neg_2 ^ x_16;
  assign px_2_18 = be_neg_2 ^ x_17;
  assign px_2_19 = be_neg_2 ^ x_18;
  assign px_2_2 = be_neg_2 ^ x_1;
  assign px_2_20 = be_neg_2 ^ x_19;
  assign px_2_21 = be_neg_2 ^ x_20;
  assign px_2_22 = be_neg_2 ^ x_21;
  assign px_2_23 = be_neg_2 ^ x_22;
  assign px_2_24 = be_neg_2 ^ x_23;
  assign px_2_25 = be_neg_2 ^ x_24;
  assign px_2_26 = be_neg_2 ^ x_25;
  assign px_2_27 = be_neg_2 ^ x_26;
  assign px_2_28 = be_neg_2 ^ x_27;
  assign px_2_29 = be_neg_2 ^ x_28;
  assign px_2_3 = be_neg_2 ^ x_2;
  assign px_2_30 = be_neg_2 ^ x_29;
  assign px_2_31 = be_neg_2 ^ x_30;
  assign px_2_32 = be_neg_2 ^ x_31;
  assign px_2_33 = be_neg_2 ^ zero;
  assign px_2_34 = be_neg_2 ^ zero;
  assign px_2_4 = be_neg_2 ^ x_3;
  assign px_2_5 = be_neg_2 ^ x_4;
  assign px_2_6 = be_neg_2 ^ x_5;
  assign px_2_7 = be_neg_2 ^ x_6;
  assign px_2_8 = be_neg_2 ^ x_7;
  assign px_2_9 = be_neg_2 ^ x_8;
  assign px_3_0 = be_neg_3;
  assign px_3_1 = be_neg_3 ^ x_0;
  assign px_3_10 = be_neg_3 ^ x_9;
  assign px_3_11 = be_neg_3 ^ x_10;
  assign px_3_12 = be_neg_3 ^ x_11;
  assign px_3_13 = be_neg_3 ^ x_12;
  assign px_3_14 = be_neg_3 ^ x_13;
  assign px_3_15 = be_neg_3 ^ x_14;
  assign px_3_16 = be_neg_3 ^ x_15;
  assign px_3_17 = be_neg_3 ^ x_16;
  assign px_3_18 = be_neg_3 ^ x_17;
  assign px_3_19 = be_neg_3 ^ x_18;
  assign px_3_2 = be_neg_3 ^ x_1;
  assign px_3_20 = be_neg_3 ^ x_19;
  assign px_3_21 = be_neg_3 ^ x_20;
  assign px_3_22 = be_neg_3 ^ x_21;
  assign px_3_23 = be_neg_3 ^ x_22;
  assign px_3_24 = be_neg_3 ^ x_23;
  assign px_3_25 = be_neg_3 ^ x_24;
  assign px_3_26 = be_neg_3 ^ x_25;
  assign px_3_27 = be_neg_3 ^ x_26;
  assign px_3_28 = be_neg_3 ^ x_27;
  assign px_3_29 = be_neg_3 ^ x_28;
  assign px_3_3 = be_neg_3 ^ x_2;
  assign px_3_30 = be_neg_3 ^ x_29;
  assign px_3_31 = be_neg_3 ^ x_30;
  assign px_3_32 = be_neg_3 ^ x_31;
  assign px_3_33 = be_neg_3 ^ zero;
  assign px_3_34 = be_neg_3 ^ zero;
  assign px_3_4 = be_neg_3 ^ x_3;
  assign px_3_5 = be_neg_3 ^ x_4;
  assign px_3_6 = be_neg_3 ^ x_5;
  assign px_3_7 = be_neg_3 ^ x_6;
  assign px_3_8 = be_neg_3 ^ x_7;
  assign px_3_9 = be_neg_3 ^ x_8;
  assign px_4_0 = be_neg_4;
  assign px_4_1 = be_neg_4 ^ x_0;
  assign px_4_10 = be_neg_4 ^ x_9;
  assign px_4_11 = be_neg_4 ^ x_10;
  assign px_4_12 = be_neg_4 ^ x_11;
  assign px_4_13 = be_neg_4 ^ x_12;
  assign px_4_14 = be_neg_4 ^ x_13;
  assign px_4_15 = be_neg_4 ^ x_14;
  assign px_4_16 = be_neg_4 ^ x_15;
  assign px_4_17 = be_neg_4 ^ x_16;
  assign px_4_18 = be_neg_4 ^ x_17;
  assign px_4_19 = be_neg_4 ^ x_18;
  assign px_4_2 = be_neg_4 ^ x_1;
  assign px_4_20 = be_neg_4 ^ x_19;
  assign px_4_21 = be_neg_4 ^ x_20;
  assign px_4_22 = be_neg_4 ^ x_21;
  assign px_4_23 = be_neg_4 ^ x_22;
  assign px_4_24 = be_neg_4 ^ x_23;
  assign px_4_25 = be_neg_4 ^ x_24;
  assign px_4_26 = be_neg_4 ^ x_25;
  assign px_4_27 = be_neg_4 ^ x_26;
  assign px_4_28 = be_neg_4 ^ x_27;
  assign px_4_29 = be_neg_4 ^ x_28;
  assign px_4_3 = be_neg_4 ^ x_2;
  assign px_4_30 = be_neg_4 ^ x_29;
  assign px_4_31 = be_neg_4 ^ x_30;
  assign px_4_32 = be_neg_4 ^ x_31;
  assign px_4_33 = be_neg_4 ^ zero;
  assign px_4_34 = be_neg_4 ^ zero;
  assign px_4_4 = be_neg_4 ^ x_3;
  assign px_4_5 = be_neg_4 ^ x_4;
  assign px_4_6 = be_neg_4 ^ x_5;
  assign px_4_7 = be_neg_4 ^ x_6;
  assign px_4_8 = be_neg_4 ^ x_7;
  assign px_4_9 = be_neg_4 ^ x_8;
  assign px_5_0 = be_neg_5;
  assign px_5_1 = be_neg_5 ^ x_0;
  assign px_5_10 = be_neg_5 ^ x_9;
  assign px_5_11 = be_neg_5 ^ x_10;
  assign px_5_12 = be_neg_5 ^ x_11;
  assign px_5_13 = be_neg_5 ^ x_12;
  assign px_5_14 = be_neg_5 ^ x_13;
  assign px_5_15 = be_neg_5 ^ x_14;
  assign px_5_16 = be_neg_5 ^ x_15;
  assign px_5_17 = be_neg_5 ^ x_16;
  assign px_5_18 = be_neg_5 ^ x_17;
  assign px_5_19 = be_neg_5 ^ x_18;
  assign px_5_2 = be_neg_5 ^ x_1;
  assign px_5_20 = be_neg_5 ^ x_19;
  assign px_5_21 = be_neg_5 ^ x_20;
  assign px_5_22 = be_neg_5 ^ x_21;
  assign px_5_23 = be_neg_5 ^ x_22;
  assign px_5_24 = be_neg_5 ^ x_23;
  assign px_5_25 = be_neg_5 ^ x_24;
  assign px_5_26 = be_neg_5 ^ x_25;
  assign px_5_27 = be_neg_5 ^ x_26;
  assign px_5_28 = be_neg_5 ^ x_27;
  assign px_5_29 = be_neg_5 ^ x_28;
  assign px_5_3 = be_neg_5 ^ x_2;
  assign px_5_30 = be_neg_5 ^ x_29;
  assign px_5_31 = be_neg_5 ^ x_30;
  assign px_5_32 = be_neg_5 ^ x_31;
  assign px_5_33 = be_neg_5 ^ zero;
  assign px_5_34 = be_neg_5 ^ zero;
  assign px_5_4 = be_neg_5 ^ x_3;
  assign px_5_5 = be_neg_5 ^ x_4;
  assign px_5_6 = be_neg_5 ^ x_5;
  assign px_5_7 = be_neg_5 ^ x_6;
  assign px_5_8 = be_neg_5 ^ x_7;
  assign px_5_9 = be_neg_5 ^ x_8;
  assign px_6_0 = be_neg_6;
  assign px_6_1 = be_neg_6 ^ x_0;
  assign px_6_10 = be_neg_6 ^ x_9;
  assign px_6_11 = be_neg_6 ^ x_10;
  assign px_6_12 = be_neg_6 ^ x_11;
  assign px_6_13 = be_neg_6 ^ x_12;
  assign px_6_14 = be_neg_6 ^ x_13;
  assign px_6_15 = be_neg_6 ^ x_14;
  assign px_6_16 = be_neg_6 ^ x_15;
  assign px_6_17 = be_neg_6 ^ x_16;
  assign px_6_18 = be_neg_6 ^ x_17;
  assign px_6_19 = be_neg_6 ^ x_18;
  assign px_6_2 = be_neg_6 ^ x_1;
  assign px_6_20 = be_neg_6 ^ x_19;
  assign px_6_21 = be_neg_6 ^ x_20;
  assign px_6_22 = be_neg_6 ^ x_21;
  assign px_6_23 = be_neg_6 ^ x_22;
  assign px_6_24 = be_neg_6 ^ x_23;
  assign px_6_25 = be_neg_6 ^ x_24;
  assign px_6_26 = be_neg_6 ^ x_25;
  assign px_6_27 = be_neg_6 ^ x_26;
  assign px_6_28 = be_neg_6 ^ x_27;
  assign px_6_29 = be_neg_6 ^ x_28;
  assign px_6_3 = be_neg_6 ^ x_2;
  assign px_6_30 = be_neg_6 ^ x_29;
  assign px_6_31 = be_neg_6 ^ x_30;
  assign px_6_32 = be_neg_6 ^ x_31;
  assign px_6_33 = be_neg_6 ^ zero;
  assign px_6_34 = be_neg_6 ^ zero;
  assign px_6_4 = be_neg_6 ^ x_3;
  assign px_6_5 = be_neg_6 ^ x_4;
  assign px_6_6 = be_neg_6 ^ x_5;
  assign px_6_7 = be_neg_6 ^ x_6;
  assign px_6_8 = be_neg_6 ^ x_7;
  assign px_6_9 = be_neg_6 ^ x_8;
  assign px_7_0 = be_neg_7;
  assign px_7_1 = be_neg_7 ^ x_0;
  assign px_7_10 = be_neg_7 ^ x_9;
  assign px_7_11 = be_neg_7 ^ x_10;
  assign px_7_12 = be_neg_7 ^ x_11;
  assign px_7_13 = be_neg_7 ^ x_12;
  assign px_7_14 = be_neg_7 ^ x_13;
  assign px_7_15 = be_neg_7 ^ x_14;
  assign px_7_16 = be_neg_7 ^ x_15;
  assign px_7_17 = be_neg_7 ^ x_16;
  assign px_7_18 = be_neg_7 ^ x_17;
  assign px_7_19 = be_neg_7 ^ x_18;
  assign px_7_2 = be_neg_7 ^ x_1;
  assign px_7_20 = be_neg_7 ^ x_19;
  assign px_7_21 = be_neg_7 ^ x_20;
  assign px_7_22 = be_neg_7 ^ x_21;
  assign px_7_23 = be_neg_7 ^ x_22;
  assign px_7_24 = be_neg_7 ^ x_23;
  assign px_7_25 = be_neg_7 ^ x_24;
  assign px_7_26 = be_neg_7 ^ x_25;
  assign px_7_27 = be_neg_7 ^ x_26;
  assign px_7_28 = be_neg_7 ^ x_27;
  assign px_7_29 = be_neg_7 ^ x_28;
  assign px_7_3 = be_neg_7 ^ x_2;
  assign px_7_30 = be_neg_7 ^ x_29;
  assign px_7_31 = be_neg_7 ^ x_30;
  assign px_7_32 = be_neg_7 ^ x_31;
  assign px_7_33 = be_neg_7 ^ zero;
  assign px_7_34 = be_neg_7 ^ zero;
  assign px_7_4 = be_neg_7 ^ x_3;
  assign px_7_5 = be_neg_7 ^ x_4;
  assign px_7_6 = be_neg_7 ^ x_5;
  assign px_7_7 = be_neg_7 ^ x_6;
  assign px_7_8 = be_neg_7 ^ x_7;
  assign px_7_9 = be_neg_7 ^ x_8;
  assign px_8_0 = be_neg_8;
  assign px_8_1 = be_neg_8 ^ x_0;
  assign px_8_10 = be_neg_8 ^ x_9;
  assign px_8_11 = be_neg_8 ^ x_10;
  assign px_8_12 = be_neg_8 ^ x_11;
  assign px_8_13 = be_neg_8 ^ x_12;
  assign px_8_14 = be_neg_8 ^ x_13;
  assign px_8_15 = be_neg_8 ^ x_14;
  assign px_8_16 = be_neg_8 ^ x_15;
  assign px_8_17 = be_neg_8 ^ x_16;
  assign px_8_18 = be_neg_8 ^ x_17;
  assign px_8_19 = be_neg_8 ^ x_18;
  assign px_8_2 = be_neg_8 ^ x_1;
  assign px_8_20 = be_neg_8 ^ x_19;
  assign px_8_21 = be_neg_8 ^ x_20;
  assign px_8_22 = be_neg_8 ^ x_21;
  assign px_8_23 = be_neg_8 ^ x_22;
  assign px_8_24 = be_neg_8 ^ x_23;
  assign px_8_25 = be_neg_8 ^ x_24;
  assign px_8_26 = be_neg_8 ^ x_25;
  assign px_8_27 = be_neg_8 ^ x_26;
  assign px_8_28 = be_neg_8 ^ x_27;
  assign px_8_29 = be_neg_8 ^ x_28;
  assign px_8_3 = be_neg_8 ^ x_2;
  assign px_8_30 = be_neg_8 ^ x_29;
  assign px_8_31 = be_neg_8 ^ x_30;
  assign px_8_32 = be_neg_8 ^ x_31;
  assign px_8_33 = be_neg_8 ^ zero;
  assign px_8_34 = be_neg_8 ^ zero;
  assign px_8_4 = be_neg_8 ^ x_3;
  assign px_8_5 = be_neg_8 ^ x_4;
  assign px_8_6 = be_neg_8 ^ x_5;
  assign px_8_7 = be_neg_8 ^ x_6;
  assign px_8_8 = be_neg_8 ^ x_7;
  assign px_8_9 = be_neg_8 ^ x_8;
  assign px_9_0 = be_neg_9;
  assign px_9_1 = be_neg_9 ^ x_0;
  assign px_9_10 = be_neg_9 ^ x_9;
  assign px_9_11 = be_neg_9 ^ x_10;
  assign px_9_12 = be_neg_9 ^ x_11;
  assign px_9_13 = be_neg_9 ^ x_12;
  assign px_9_14 = be_neg_9 ^ x_13;
  assign px_9_15 = be_neg_9 ^ x_14;
  assign px_9_16 = be_neg_9 ^ x_15;
  assign px_9_17 = be_neg_9 ^ x_16;
  assign px_9_18 = be_neg_9 ^ x_17;
  assign px_9_19 = be_neg_9 ^ x_18;
  assign px_9_2 = be_neg_9 ^ x_1;
  assign px_9_20 = be_neg_9 ^ x_19;
  assign px_9_21 = be_neg_9 ^ x_20;
  assign px_9_22 = be_neg_9 ^ x_21;
  assign px_9_23 = be_neg_9 ^ x_22;
  assign px_9_24 = be_neg_9 ^ x_23;
  assign px_9_25 = be_neg_9 ^ x_24;
  assign px_9_26 = be_neg_9 ^ x_25;
  assign px_9_27 = be_neg_9 ^ x_26;
  assign px_9_28 = be_neg_9 ^ x_27;
  assign px_9_29 = be_neg_9 ^ x_28;
  assign px_9_3 = be_neg_9 ^ x_2;
  assign px_9_30 = be_neg_9 ^ x_29;
  assign px_9_31 = be_neg_9 ^ x_30;
  assign px_9_32 = be_neg_9 ^ x_31;
  assign px_9_33 = be_neg_9 ^ zero;
  assign px_9_34 = be_neg_9 ^ zero;
  assign px_9_4 = be_neg_9 ^ x_3;
  assign px_9_5 = be_neg_9 ^ x_4;
  assign px_9_6 = be_neg_9 ^ x_5;
  assign px_9_7 = be_neg_9 ^ x_6;
  assign px_9_8 = be_neg_9 ^ x_7;
  assign px_9_9 = be_neg_9 ^ x_8;
  assign x_0 = multiplicand[0];
  assign x_1 = multiplicand[1];
  assign x_10 = multiplicand[10];
  assign x_11 = multiplicand[11];
  assign x_12 = multiplicand[12];
  assign x_13 = multiplicand[13];
  assign x_14 = multiplicand[14];
  assign x_15 = multiplicand[15];
  assign x_16 = multiplicand[16];
  assign x_17 = multiplicand[17];
  assign x_18 = multiplicand[18];
  assign x_19 = multiplicand[19];
  assign x_2 = multiplicand[2];
  assign x_20 = multiplicand[20];
  assign x_21 = multiplicand[21];
  assign x_22 = multiplicand[22];
  assign x_23 = multiplicand[23];
  assign x_24 = multiplicand[24];
  assign x_25 = multiplicand[25];
  assign x_26 = multiplicand[26];
  assign x_27 = multiplicand[27];
  assign x_28 = multiplicand[28];
  assign x_29 = multiplicand[29];
  assign x_3 = multiplicand[3];
  assign x_30 = multiplicand[30];
  assign x_31 = multiplicand[31];
  assign x_4 = multiplicand[4];
  assign x_5 = multiplicand[5];
  assign x_6 = multiplicand[6];
  assign x_7 = multiplicand[7];
  assign x_8 = multiplicand[8];
  assign x_9 = multiplicand[9];
  assign y_0 = multiplier[0];
  assign y_1 = multiplier[1];
  assign y_10 = multiplier[10];
  assign y_11 = multiplier[11];
  assign y_12 = multiplier[12];
  assign y_13 = multiplier[13];
  assign y_14 = multiplier[14];
  assign y_15 = multiplier[15];
  assign y_16 = multiplier[16];
  assign y_17 = multiplier[17];
  assign y_18 = multiplier[18];
  assign y_19 = multiplier[19];
  assign y_2 = multiplier[2];
  assign y_20 = multiplier[20];
  assign y_21 = multiplier[21];
  assign y_22 = multiplier[22];
  assign y_23 = multiplier[23];
  assign y_24 = multiplier[24];
  assign y_25 = multiplier[25];
  assign y_26 = multiplier[26];
  assign y_27 = multiplier[27];
  assign y_28 = multiplier[28];
  assign y_29 = multiplier[29];
  assign y_3 = multiplier[3];
  assign y_30 = multiplier[30];
  assign y_31 = multiplier[31];
  assign y_4 = multiplier[4];
  assign y_5 = multiplier[5];
  assign y_6 = multiplier[6];
  assign y_7 = multiplier[7];
  assign y_8 = multiplier[8];
  assign y_9 = multiplier[9];
  assign zero = 1'b0;
  wire pp_0_0_0;
  wire pp_0_0_1;
  wire pp_0_1_0;
  wire pp_0_2_0;
  wire pp_0_2_1;
  wire pp_0_2_2;
  wire pp_0_3_0;
  wire pp_0_3_1;
  wire pp_0_4_0;
  wire pp_0_4_1;
  wire pp_0_4_2;
  wire pp_0_4_3;
  wire pp_0_5_0;
  wire pp_0_5_1;
  wire pp_0_5_2;
  wire pp_0_6_0;
  wire pp_0_6_1;
  wire pp_0_6_2;
  wire pp_0_6_3;
  wire pp_0_6_4;
  wire pp_0_7_0;
  wire pp_0_7_1;
  wire pp_0_7_2;
  wire pp_0_7_3;
  wire pp_0_8_0;
  wire pp_0_8_1;
  wire pp_0_8_2;
  wire pp_0_8_3;
  wire pp_0_8_4;
  wire pp_0_8_5;
  wire pp_0_9_0;
  wire pp_0_9_1;
  wire pp_0_9_2;
  wire pp_0_9_3;
  wire pp_0_9_4;
  wire pp_0_10_0;
  wire pp_0_10_1;
  wire pp_0_10_2;
  wire pp_0_10_3;
  wire pp_0_10_4;
  wire pp_0_10_5;
  wire pp_0_10_6;
  wire pp_0_11_0;
  wire pp_0_11_1;
  wire pp_0_11_2;
  wire pp_0_11_3;
  wire pp_0_11_4;
  wire pp_0_11_5;
  wire pp_0_12_0;
  wire pp_0_12_1;
  wire pp_0_12_2;
  wire pp_0_12_3;
  wire pp_0_12_4;
  wire pp_0_12_5;
  wire pp_0_12_6;
  wire pp_0_12_7;
  wire pp_0_13_0;
  wire pp_0_13_1;
  wire pp_0_13_2;
  wire pp_0_13_3;
  wire pp_0_13_4;
  wire pp_0_13_5;
  wire pp_0_13_6;
  wire pp_0_14_0;
  wire pp_0_14_1;
  wire pp_0_14_2;
  wire pp_0_14_3;
  wire pp_0_14_4;
  wire pp_0_14_5;
  wire pp_0_14_6;
  wire pp_0_14_7;
  wire pp_0_14_8;
  wire pp_0_15_0;
  wire pp_0_15_1;
  wire pp_0_15_2;
  wire pp_0_15_3;
  wire pp_0_15_4;
  wire pp_0_15_5;
  wire pp_0_15_6;
  wire pp_0_15_7;
  wire pp_0_16_0;
  wire pp_0_16_1;
  wire pp_0_16_2;
  wire pp_0_16_3;
  wire pp_0_16_4;
  wire pp_0_16_5;
  wire pp_0_16_6;
  wire pp_0_16_7;
  wire pp_0_16_8;
  wire pp_0_16_9;
  wire pp_0_17_0;
  wire pp_0_17_1;
  wire pp_0_17_2;
  wire pp_0_17_3;
  wire pp_0_17_4;
  wire pp_0_17_5;
  wire pp_0_17_6;
  wire pp_0_17_7;
  wire pp_0_17_8;
  wire pp_0_18_0;
  wire pp_0_18_1;
  wire pp_0_18_2;
  wire pp_0_18_3;
  wire pp_0_18_4;
  wire pp_0_18_5;
  wire pp_0_18_6;
  wire pp_0_18_7;
  wire pp_0_18_8;
  wire pp_0_18_9;
  wire pp_0_18_10;
  wire pp_0_19_0;
  wire pp_0_19_1;
  wire pp_0_19_2;
  wire pp_0_19_3;
  wire pp_0_19_4;
  wire pp_0_19_5;
  wire pp_0_19_6;
  wire pp_0_19_7;
  wire pp_0_19_8;
  wire pp_0_19_9;
  wire pp_0_20_0;
  wire pp_0_20_1;
  wire pp_0_20_2;
  wire pp_0_20_3;
  wire pp_0_20_4;
  wire pp_0_20_5;
  wire pp_0_20_6;
  wire pp_0_20_7;
  wire pp_0_20_8;
  wire pp_0_20_9;
  wire pp_0_20_10;
  wire pp_0_20_11;
  wire pp_0_21_0;
  wire pp_0_21_1;
  wire pp_0_21_2;
  wire pp_0_21_3;
  wire pp_0_21_4;
  wire pp_0_21_5;
  wire pp_0_21_6;
  wire pp_0_21_7;
  wire pp_0_21_8;
  wire pp_0_21_9;
  wire pp_0_21_10;
  wire pp_0_22_0;
  wire pp_0_22_1;
  wire pp_0_22_2;
  wire pp_0_22_3;
  wire pp_0_22_4;
  wire pp_0_22_5;
  wire pp_0_22_6;
  wire pp_0_22_7;
  wire pp_0_22_8;
  wire pp_0_22_9;
  wire pp_0_22_10;
  wire pp_0_22_11;
  wire pp_0_22_12;
  wire pp_0_23_0;
  wire pp_0_23_1;
  wire pp_0_23_2;
  wire pp_0_23_3;
  wire pp_0_23_4;
  wire pp_0_23_5;
  wire pp_0_23_6;
  wire pp_0_23_7;
  wire pp_0_23_8;
  wire pp_0_23_9;
  wire pp_0_23_10;
  wire pp_0_23_11;
  wire pp_0_24_0;
  wire pp_0_24_1;
  wire pp_0_24_2;
  wire pp_0_24_3;
  wire pp_0_24_4;
  wire pp_0_24_5;
  wire pp_0_24_6;
  wire pp_0_24_7;
  wire pp_0_24_8;
  wire pp_0_24_9;
  wire pp_0_24_10;
  wire pp_0_24_11;
  wire pp_0_24_12;
  wire pp_0_24_13;
  wire pp_0_25_0;
  wire pp_0_25_1;
  wire pp_0_25_2;
  wire pp_0_25_3;
  wire pp_0_25_4;
  wire pp_0_25_5;
  wire pp_0_25_6;
  wire pp_0_25_7;
  wire pp_0_25_8;
  wire pp_0_25_9;
  wire pp_0_25_10;
  wire pp_0_25_11;
  wire pp_0_25_12;
  wire pp_0_26_0;
  wire pp_0_26_1;
  wire pp_0_26_2;
  wire pp_0_26_3;
  wire pp_0_26_4;
  wire pp_0_26_5;
  wire pp_0_26_6;
  wire pp_0_26_7;
  wire pp_0_26_8;
  wire pp_0_26_9;
  wire pp_0_26_10;
  wire pp_0_26_11;
  wire pp_0_26_12;
  wire pp_0_26_13;
  wire pp_0_26_14;
  wire pp_0_27_0;
  wire pp_0_27_1;
  wire pp_0_27_2;
  wire pp_0_27_3;
  wire pp_0_27_4;
  wire pp_0_27_5;
  wire pp_0_27_6;
  wire pp_0_27_7;
  wire pp_0_27_8;
  wire pp_0_27_9;
  wire pp_0_27_10;
  wire pp_0_27_11;
  wire pp_0_27_12;
  wire pp_0_27_13;
  wire pp_0_28_0;
  wire pp_0_28_1;
  wire pp_0_28_2;
  wire pp_0_28_3;
  wire pp_0_28_4;
  wire pp_0_28_5;
  wire pp_0_28_6;
  wire pp_0_28_7;
  wire pp_0_28_8;
  wire pp_0_28_9;
  wire pp_0_28_10;
  wire pp_0_28_11;
  wire pp_0_28_12;
  wire pp_0_28_13;
  wire pp_0_28_14;
  wire pp_0_28_15;
  wire pp_0_29_0;
  wire pp_0_29_1;
  wire pp_0_29_2;
  wire pp_0_29_3;
  wire pp_0_29_4;
  wire pp_0_29_5;
  wire pp_0_29_6;
  wire pp_0_29_7;
  wire pp_0_29_8;
  wire pp_0_29_9;
  wire pp_0_29_10;
  wire pp_0_29_11;
  wire pp_0_29_12;
  wire pp_0_29_13;
  wire pp_0_29_14;
  wire pp_0_30_0;
  wire pp_0_30_1;
  wire pp_0_30_2;
  wire pp_0_30_3;
  wire pp_0_30_4;
  wire pp_0_30_5;
  wire pp_0_30_6;
  wire pp_0_30_7;
  wire pp_0_30_8;
  wire pp_0_30_9;
  wire pp_0_30_10;
  wire pp_0_30_11;
  wire pp_0_30_12;
  wire pp_0_30_13;
  wire pp_0_30_14;
  wire pp_0_30_15;
  wire pp_0_30_16;
  wire pp_0_31_0;
  wire pp_0_31_1;
  wire pp_0_31_2;
  wire pp_0_31_3;
  wire pp_0_31_4;
  wire pp_0_31_5;
  wire pp_0_31_6;
  wire pp_0_31_7;
  wire pp_0_31_8;
  wire pp_0_31_9;
  wire pp_0_31_10;
  wire pp_0_31_11;
  wire pp_0_31_12;
  wire pp_0_31_13;
  wire pp_0_31_14;
  wire pp_0_31_15;
  wire pp_0_32_0;
  wire pp_0_32_1;
  wire pp_0_32_2;
  wire pp_0_32_3;
  wire pp_0_32_4;
  wire pp_0_32_5;
  wire pp_0_32_6;
  wire pp_0_32_7;
  wire pp_0_32_8;
  wire pp_0_32_9;
  wire pp_0_32_10;
  wire pp_0_32_11;
  wire pp_0_32_12;
  wire pp_0_32_13;
  wire pp_0_32_14;
  wire pp_0_32_15;
  wire pp_0_32_16;
  wire pp_0_33_0;
  wire pp_0_33_1;
  wire pp_0_33_2;
  wire pp_0_33_3;
  wire pp_0_33_4;
  wire pp_0_33_5;
  wire pp_0_33_6;
  wire pp_0_33_7;
  wire pp_0_33_8;
  wire pp_0_33_9;
  wire pp_0_33_10;
  wire pp_0_33_11;
  wire pp_0_33_12;
  wire pp_0_33_13;
  wire pp_0_33_14;
  wire pp_0_33_15;
  wire pp_0_33_16;
  wire pp_0_34_0;
  wire pp_0_34_1;
  wire pp_0_34_2;
  wire pp_0_34_3;
  wire pp_0_34_4;
  wire pp_0_34_5;
  wire pp_0_34_6;
  wire pp_0_34_7;
  wire pp_0_34_8;
  wire pp_0_34_9;
  wire pp_0_34_10;
  wire pp_0_34_11;
  wire pp_0_34_12;
  wire pp_0_34_13;
  wire pp_0_34_14;
  wire pp_0_34_15;
  wire pp_0_34_16;
  wire pp_0_35_0;
  wire pp_0_35_1;
  wire pp_0_35_2;
  wire pp_0_35_3;
  wire pp_0_35_4;
  wire pp_0_35_5;
  wire pp_0_35_6;
  wire pp_0_35_7;
  wire pp_0_35_8;
  wire pp_0_35_9;
  wire pp_0_35_10;
  wire pp_0_35_11;
  wire pp_0_35_12;
  wire pp_0_35_13;
  wire pp_0_35_14;
  wire pp_0_35_15;
  wire pp_0_35_16;
  wire pp_0_36_0;
  wire pp_0_36_1;
  wire pp_0_36_2;
  wire pp_0_36_3;
  wire pp_0_36_4;
  wire pp_0_36_5;
  wire pp_0_36_6;
  wire pp_0_36_7;
  wire pp_0_36_8;
  wire pp_0_36_9;
  wire pp_0_36_10;
  wire pp_0_36_11;
  wire pp_0_36_12;
  wire pp_0_36_13;
  wire pp_0_36_14;
  wire pp_0_36_15;
  wire pp_0_37_0;
  wire pp_0_37_1;
  wire pp_0_37_2;
  wire pp_0_37_3;
  wire pp_0_37_4;
  wire pp_0_37_5;
  wire pp_0_37_6;
  wire pp_0_37_7;
  wire pp_0_37_8;
  wire pp_0_37_9;
  wire pp_0_37_10;
  wire pp_0_37_11;
  wire pp_0_37_12;
  wire pp_0_37_13;
  wire pp_0_37_14;
  wire pp_0_38_0;
  wire pp_0_38_1;
  wire pp_0_38_2;
  wire pp_0_38_3;
  wire pp_0_38_4;
  wire pp_0_38_5;
  wire pp_0_38_6;
  wire pp_0_38_7;
  wire pp_0_38_8;
  wire pp_0_38_9;
  wire pp_0_38_10;
  wire pp_0_38_11;
  wire pp_0_38_12;
  wire pp_0_38_13;
  wire pp_0_38_14;
  wire pp_0_39_0;
  wire pp_0_39_1;
  wire pp_0_39_2;
  wire pp_0_39_3;
  wire pp_0_39_4;
  wire pp_0_39_5;
  wire pp_0_39_6;
  wire pp_0_39_7;
  wire pp_0_39_8;
  wire pp_0_39_9;
  wire pp_0_39_10;
  wire pp_0_39_11;
  wire pp_0_39_12;
  wire pp_0_39_13;
  wire pp_0_40_0;
  wire pp_0_40_1;
  wire pp_0_40_2;
  wire pp_0_40_3;
  wire pp_0_40_4;
  wire pp_0_40_5;
  wire pp_0_40_6;
  wire pp_0_40_7;
  wire pp_0_40_8;
  wire pp_0_40_9;
  wire pp_0_40_10;
  wire pp_0_40_11;
  wire pp_0_40_12;
  wire pp_0_40_13;
  wire pp_0_41_0;
  wire pp_0_41_1;
  wire pp_0_41_2;
  wire pp_0_41_3;
  wire pp_0_41_4;
  wire pp_0_41_5;
  wire pp_0_41_6;
  wire pp_0_41_7;
  wire pp_0_41_8;
  wire pp_0_41_9;
  wire pp_0_41_10;
  wire pp_0_41_11;
  wire pp_0_41_12;
  wire pp_0_42_0;
  wire pp_0_42_1;
  wire pp_0_42_2;
  wire pp_0_42_3;
  wire pp_0_42_4;
  wire pp_0_42_5;
  wire pp_0_42_6;
  wire pp_0_42_7;
  wire pp_0_42_8;
  wire pp_0_42_9;
  wire pp_0_42_10;
  wire pp_0_42_11;
  wire pp_0_42_12;
  wire pp_0_43_0;
  wire pp_0_43_1;
  wire pp_0_43_2;
  wire pp_0_43_3;
  wire pp_0_43_4;
  wire pp_0_43_5;
  wire pp_0_43_6;
  wire pp_0_43_7;
  wire pp_0_43_8;
  wire pp_0_43_9;
  wire pp_0_43_10;
  wire pp_0_43_11;
  wire pp_0_44_0;
  wire pp_0_44_1;
  wire pp_0_44_2;
  wire pp_0_44_3;
  wire pp_0_44_4;
  wire pp_0_44_5;
  wire pp_0_44_6;
  wire pp_0_44_7;
  wire pp_0_44_8;
  wire pp_0_44_9;
  wire pp_0_44_10;
  wire pp_0_44_11;
  wire pp_0_45_0;
  wire pp_0_45_1;
  wire pp_0_45_2;
  wire pp_0_45_3;
  wire pp_0_45_4;
  wire pp_0_45_5;
  wire pp_0_45_6;
  wire pp_0_45_7;
  wire pp_0_45_8;
  wire pp_0_45_9;
  wire pp_0_45_10;
  wire pp_0_46_0;
  wire pp_0_46_1;
  wire pp_0_46_2;
  wire pp_0_46_3;
  wire pp_0_46_4;
  wire pp_0_46_5;
  wire pp_0_46_6;
  wire pp_0_46_7;
  wire pp_0_46_8;
  wire pp_0_46_9;
  wire pp_0_46_10;
  wire pp_0_47_0;
  wire pp_0_47_1;
  wire pp_0_47_2;
  wire pp_0_47_3;
  wire pp_0_47_4;
  wire pp_0_47_5;
  wire pp_0_47_6;
  wire pp_0_47_7;
  wire pp_0_47_8;
  wire pp_0_47_9;
  wire pp_0_48_0;
  wire pp_0_48_1;
  wire pp_0_48_2;
  wire pp_0_48_3;
  wire pp_0_48_4;
  wire pp_0_48_5;
  wire pp_0_48_6;
  wire pp_0_48_7;
  wire pp_0_48_8;
  wire pp_0_48_9;
  wire pp_0_49_0;
  wire pp_0_49_1;
  wire pp_0_49_2;
  wire pp_0_49_3;
  wire pp_0_49_4;
  wire pp_0_49_5;
  wire pp_0_49_6;
  wire pp_0_49_7;
  wire pp_0_49_8;
  wire pp_0_50_0;
  wire pp_0_50_1;
  wire pp_0_50_2;
  wire pp_0_50_3;
  wire pp_0_50_4;
  wire pp_0_50_5;
  wire pp_0_50_6;
  wire pp_0_50_7;
  wire pp_0_50_8;
  wire pp_0_51_0;
  wire pp_0_51_1;
  wire pp_0_51_2;
  wire pp_0_51_3;
  wire pp_0_51_4;
  wire pp_0_51_5;
  wire pp_0_51_6;
  wire pp_0_51_7;
  wire pp_0_52_0;
  wire pp_0_52_1;
  wire pp_0_52_2;
  wire pp_0_52_3;
  wire pp_0_52_4;
  wire pp_0_52_5;
  wire pp_0_52_6;
  wire pp_0_52_7;
  wire pp_0_53_0;
  wire pp_0_53_1;
  wire pp_0_53_2;
  wire pp_0_53_3;
  wire pp_0_53_4;
  wire pp_0_53_5;
  wire pp_0_53_6;
  wire pp_0_54_0;
  wire pp_0_54_1;
  wire pp_0_54_2;
  wire pp_0_54_3;
  wire pp_0_54_4;
  wire pp_0_54_5;
  wire pp_0_54_6;
  wire pp_0_55_0;
  wire pp_0_55_1;
  wire pp_0_55_2;
  wire pp_0_55_3;
  wire pp_0_55_4;
  wire pp_0_55_5;
  wire pp_0_56_0;
  wire pp_0_56_1;
  wire pp_0_56_2;
  wire pp_0_56_3;
  wire pp_0_56_4;
  wire pp_0_56_5;
  wire pp_0_57_0;
  wire pp_0_57_1;
  wire pp_0_57_2;
  wire pp_0_57_3;
  wire pp_0_57_4;
  wire pp_0_58_0;
  wire pp_0_58_1;
  wire pp_0_58_2;
  wire pp_0_58_3;
  wire pp_0_58_4;
  wire pp_0_59_0;
  wire pp_0_59_1;
  wire pp_0_59_2;
  wire pp_0_59_3;
  wire pp_0_60_0;
  wire pp_0_60_1;
  wire pp_0_60_2;
  wire pp_0_60_3;
  wire pp_0_61_0;
  wire pp_0_61_1;
  wire pp_0_61_2;
  wire pp_0_62_0;
  wire pp_0_62_1;
  wire pp_0_62_2;
  wire pp_0_63_0;
  wire pp_0_63_1;
  wire pp_1_0_0;
  wire pp_1_0_1;
  wire pp_1_1_0;
  wire pp_1_2_0;
  wire pp_1_2_1;
  wire pp_1_3_0;
  wire pp_1_3_1;
  wire pp_1_4_0;
  wire pp_1_4_1;
  wire pp_1_4_2;
  wire pp_1_4_3;
  wire pp_1_4_4;
  wire pp_1_5_0;
  wire pp_1_5_1;
  wire pp_1_5_2;
  wire pp_1_6_0;
  wire pp_1_6_1;
  wire pp_1_6_2;
  wire pp_1_7_0;
  wire pp_1_7_1;
  wire pp_1_7_2;
  wire pp_1_8_0;
  wire pp_1_8_1;
  wire pp_1_8_2;
  wire pp_1_9_0;
  wire pp_1_9_1;
  wire pp_1_9_2;
  wire pp_1_9_3;
  wire pp_1_9_4;
  wire pp_1_9_5;
  wire pp_1_9_6;
  wire pp_1_10_0;
  wire pp_1_10_1;
  wire pp_1_10_2;
  wire pp_1_11_0;
  wire pp_1_11_1;
  wire pp_1_11_2;
  wire pp_1_11_3;
  wire pp_1_12_0;
  wire pp_1_12_1;
  wire pp_1_12_2;
  wire pp_1_12_3;
  wire pp_1_12_4;
  wire pp_1_12_5;
  wire pp_1_13_0;
  wire pp_1_13_1;
  wire pp_1_13_2;
  wire pp_1_13_3;
  wire pp_1_13_4;
  wire pp_1_13_5;
  wire pp_1_13_6;
  wire pp_1_14_0;
  wire pp_1_14_1;
  wire pp_1_14_2;
  wire pp_1_14_3;
  wire pp_1_15_0;
  wire pp_1_15_1;
  wire pp_1_15_2;
  wire pp_1_15_3;
  wire pp_1_15_4;
  wire pp_1_15_5;
  wire pp_1_15_6;
  wire pp_1_16_0;
  wire pp_1_16_1;
  wire pp_1_16_2;
  wire pp_1_16_3;
  wire pp_1_16_4;
  wire pp_1_16_5;
  wire pp_1_17_0;
  wire pp_1_17_1;
  wire pp_1_17_2;
  wire pp_1_17_3;
  wire pp_1_17_4;
  wire pp_1_17_5;
  wire pp_1_18_0;
  wire pp_1_18_1;
  wire pp_1_18_2;
  wire pp_1_18_3;
  wire pp_1_18_4;
  wire pp_1_18_5;
  wire pp_1_18_6;
  wire pp_1_18_7;
  wire pp_1_18_8;
  wire pp_1_18_9;
  wire pp_1_19_0;
  wire pp_1_19_1;
  wire pp_1_19_2;
  wire pp_1_19_3;
  wire pp_1_19_4;
  wire pp_1_19_5;
  wire pp_1_20_0;
  wire pp_1_20_1;
  wire pp_1_20_2;
  wire pp_1_20_3;
  wire pp_1_20_4;
  wire pp_1_20_5;
  wire pp_1_20_6;
  wire pp_1_21_0;
  wire pp_1_21_1;
  wire pp_1_21_2;
  wire pp_1_21_3;
  wire pp_1_21_4;
  wire pp_1_21_5;
  wire pp_1_21_6;
  wire pp_1_21_7;
  wire pp_1_21_8;
  wire pp_1_22_0;
  wire pp_1_22_1;
  wire pp_1_22_2;
  wire pp_1_22_3;
  wire pp_1_22_4;
  wire pp_1_22_5;
  wire pp_1_22_6;
  wire pp_1_22_7;
  wire pp_1_23_0;
  wire pp_1_23_1;
  wire pp_1_23_2;
  wire pp_1_23_3;
  wire pp_1_23_4;
  wire pp_1_23_5;
  wire pp_1_23_6;
  wire pp_1_23_7;
  wire pp_1_24_0;
  wire pp_1_24_1;
  wire pp_1_24_2;
  wire pp_1_24_3;
  wire pp_1_24_4;
  wire pp_1_24_5;
  wire pp_1_24_6;
  wire pp_1_24_7;
  wire pp_1_24_8;
  wire pp_1_24_9;
  wire pp_1_25_0;
  wire pp_1_25_1;
  wire pp_1_25_2;
  wire pp_1_25_3;
  wire pp_1_25_4;
  wire pp_1_25_5;
  wire pp_1_25_6;
  wire pp_1_25_7;
  wire pp_1_25_8;
  wire pp_1_26_0;
  wire pp_1_26_1;
  wire pp_1_26_2;
  wire pp_1_26_3;
  wire pp_1_26_4;
  wire pp_1_26_5;
  wire pp_1_26_6;
  wire pp_1_26_7;
  wire pp_1_26_8;
  wire pp_1_27_0;
  wire pp_1_27_1;
  wire pp_1_27_2;
  wire pp_1_27_3;
  wire pp_1_27_4;
  wire pp_1_27_5;
  wire pp_1_27_6;
  wire pp_1_27_7;
  wire pp_1_27_8;
  wire pp_1_27_9;
  wire pp_1_27_10;
  wire pp_1_27_11;
  wire pp_1_27_12;
  wire pp_1_28_0;
  wire pp_1_28_1;
  wire pp_1_28_2;
  wire pp_1_28_3;
  wire pp_1_28_4;
  wire pp_1_28_5;
  wire pp_1_28_6;
  wire pp_1_28_7;
  wire pp_1_28_8;
  wire pp_1_29_0;
  wire pp_1_29_1;
  wire pp_1_29_2;
  wire pp_1_29_3;
  wire pp_1_29_4;
  wire pp_1_29_5;
  wire pp_1_29_6;
  wire pp_1_29_7;
  wire pp_1_29_8;
  wire pp_1_29_9;
  wire pp_1_30_0;
  wire pp_1_30_1;
  wire pp_1_30_2;
  wire pp_1_30_3;
  wire pp_1_30_4;
  wire pp_1_30_5;
  wire pp_1_30_6;
  wire pp_1_30_7;
  wire pp_1_30_8;
  wire pp_1_30_9;
  wire pp_1_30_10;
  wire pp_1_30_11;
  wire pp_1_31_0;
  wire pp_1_31_1;
  wire pp_1_31_2;
  wire pp_1_31_3;
  wire pp_1_31_4;
  wire pp_1_31_5;
  wire pp_1_31_6;
  wire pp_1_31_7;
  wire pp_1_31_8;
  wire pp_1_31_9;
  wire pp_1_31_10;
  wire pp_1_31_11;
  wire pp_1_32_0;
  wire pp_1_32_1;
  wire pp_1_32_2;
  wire pp_1_32_3;
  wire pp_1_32_4;
  wire pp_1_32_5;
  wire pp_1_32_6;
  wire pp_1_32_7;
  wire pp_1_32_8;
  wire pp_1_32_9;
  wire pp_1_32_10;
  wire pp_1_32_11;
  wire pp_1_33_0;
  wire pp_1_33_1;
  wire pp_1_33_2;
  wire pp_1_33_3;
  wire pp_1_33_4;
  wire pp_1_33_5;
  wire pp_1_33_6;
  wire pp_1_33_7;
  wire pp_1_33_8;
  wire pp_1_33_9;
  wire pp_1_33_10;
  wire pp_1_33_11;
  wire pp_1_34_0;
  wire pp_1_34_1;
  wire pp_1_34_2;
  wire pp_1_34_3;
  wire pp_1_34_4;
  wire pp_1_34_5;
  wire pp_1_34_6;
  wire pp_1_34_7;
  wire pp_1_34_8;
  wire pp_1_34_9;
  wire pp_1_34_10;
  wire pp_1_34_11;
  wire pp_1_35_0;
  wire pp_1_35_1;
  wire pp_1_35_2;
  wire pp_1_35_3;
  wire pp_1_35_4;
  wire pp_1_35_5;
  wire pp_1_35_6;
  wire pp_1_35_7;
  wire pp_1_35_8;
  wire pp_1_35_9;
  wire pp_1_35_10;
  wire pp_1_35_11;
  wire pp_1_36_0;
  wire pp_1_36_1;
  wire pp_1_36_2;
  wire pp_1_36_3;
  wire pp_1_36_4;
  wire pp_1_36_5;
  wire pp_1_36_6;
  wire pp_1_36_7;
  wire pp_1_36_8;
  wire pp_1_36_9;
  wire pp_1_36_10;
  wire pp_1_37_0;
  wire pp_1_37_1;
  wire pp_1_37_2;
  wire pp_1_37_3;
  wire pp_1_37_4;
  wire pp_1_37_5;
  wire pp_1_37_6;
  wire pp_1_37_7;
  wire pp_1_37_8;
  wire pp_1_37_9;
  wire pp_1_37_10;
  wire pp_1_37_11;
  wire pp_1_38_0;
  wire pp_1_38_1;
  wire pp_1_38_2;
  wire pp_1_38_3;
  wire pp_1_38_4;
  wire pp_1_38_5;
  wire pp_1_38_6;
  wire pp_1_38_7;
  wire pp_1_38_8;
  wire pp_1_39_0;
  wire pp_1_39_1;
  wire pp_1_39_2;
  wire pp_1_39_3;
  wire pp_1_39_4;
  wire pp_1_39_5;
  wire pp_1_39_6;
  wire pp_1_39_7;
  wire pp_1_39_8;
  wire pp_1_39_9;
  wire pp_1_39_10;
  wire pp_1_40_0;
  wire pp_1_40_1;
  wire pp_1_40_2;
  wire pp_1_40_3;
  wire pp_1_40_4;
  wire pp_1_40_5;
  wire pp_1_40_6;
  wire pp_1_40_7;
  wire pp_1_40_8;
  wire pp_1_40_9;
  wire pp_1_41_0;
  wire pp_1_41_1;
  wire pp_1_41_2;
  wire pp_1_41_3;
  wire pp_1_41_4;
  wire pp_1_41_5;
  wire pp_1_41_6;
  wire pp_1_41_7;
  wire pp_1_41_8;
  wire pp_1_42_0;
  wire pp_1_42_1;
  wire pp_1_42_2;
  wire pp_1_42_3;
  wire pp_1_42_4;
  wire pp_1_42_5;
  wire pp_1_42_6;
  wire pp_1_42_7;
  wire pp_1_42_8;
  wire pp_1_43_0;
  wire pp_1_43_1;
  wire pp_1_43_2;
  wire pp_1_43_3;
  wire pp_1_43_4;
  wire pp_1_43_5;
  wire pp_1_43_6;
  wire pp_1_43_7;
  wire pp_1_43_8;
  wire pp_1_43_9;
  wire pp_1_43_10;
  wire pp_1_43_11;
  wire pp_1_44_0;
  wire pp_1_44_1;
  wire pp_1_44_2;
  wire pp_1_44_3;
  wire pp_1_44_4;
  wire pp_1_44_5;
  wire pp_1_45_0;
  wire pp_1_45_1;
  wire pp_1_45_2;
  wire pp_1_45_3;
  wire pp_1_45_4;
  wire pp_1_45_5;
  wire pp_1_45_6;
  wire pp_1_45_7;
  wire pp_1_45_8;
  wire pp_1_45_9;
  wire pp_1_45_10;
  wire pp_1_45_11;
  wire pp_1_45_12;
  wire pp_1_46_0;
  wire pp_1_46_1;
  wire pp_1_46_2;
  wire pp_1_46_3;
  wire pp_1_46_4;
  wire pp_1_46_5;
  wire pp_1_46_6;
  wire pp_1_46_7;
  wire pp_1_46_8;
  wire pp_1_47_0;
  wire pp_1_47_1;
  wire pp_1_47_2;
  wire pp_1_47_3;
  wire pp_1_47_4;
  wire pp_1_47_5;
  wire pp_1_48_0;
  wire pp_1_48_1;
  wire pp_1_48_2;
  wire pp_1_48_3;
  wire pp_1_48_4;
  wire pp_1_48_5;
  wire pp_1_48_6;
  wire pp_1_48_7;
  wire pp_1_48_8;
  wire pp_1_49_0;
  wire pp_1_49_1;
  wire pp_1_49_2;
  wire pp_1_49_3;
  wire pp_1_49_4;
  wire pp_1_50_0;
  wire pp_1_50_1;
  wire pp_1_50_2;
  wire pp_1_50_3;
  wire pp_1_50_4;
  wire pp_1_50_5;
  wire pp_1_51_0;
  wire pp_1_51_1;
  wire pp_1_51_2;
  wire pp_1_51_3;
  wire pp_1_51_4;
  wire pp_1_51_5;
  wire pp_1_51_6;
  wire pp_1_52_0;
  wire pp_1_52_1;
  wire pp_1_52_2;
  wire pp_1_52_3;
  wire pp_1_52_4;
  wire pp_1_52_5;
  wire pp_1_53_0;
  wire pp_1_53_1;
  wire pp_1_53_2;
  wire pp_1_53_3;
  wire pp_1_53_4;
  wire pp_1_53_5;
  wire pp_1_53_6;
  wire pp_1_53_7;
  wire pp_1_53_8;
  wire pp_1_54_0;
  wire pp_1_54_1;
  wire pp_1_54_2;
  wire pp_1_55_0;
  wire pp_1_55_1;
  wire pp_1_55_2;
  wire pp_1_55_3;
  wire pp_1_56_0;
  wire pp_1_56_1;
  wire pp_1_56_2;
  wire pp_1_56_3;
  wire pp_1_56_4;
  wire pp_1_56_5;
  wire pp_1_56_6;
  wire pp_1_56_7;
  wire pp_1_57_0;
  wire pp_1_57_1;
  wire pp_1_57_2;
  wire pp_1_58_0;
  wire pp_1_58_1;
  wire pp_1_58_2;
  wire pp_1_58_3;
  wire pp_1_58_4;
  wire pp_1_58_5;
  wire pp_1_59_0;
  wire pp_1_59_1;
  wire pp_1_60_0;
  wire pp_1_60_1;
  wire pp_1_60_2;
  wire pp_1_61_0;
  wire pp_1_61_1;
  wire pp_1_61_2;
  wire pp_1_61_3;
  wire pp_1_62_0;
  wire pp_1_62_1;
  wire pp_1_62_2;
  wire pp_1_63_0;
  wire pp_1_63_1;
  wire pp_2_0_0;
  wire pp_2_0_1;
  wire pp_2_1_0;
  wire pp_2_2_0;
  wire pp_2_2_1;
  wire pp_2_3_0;
  wire pp_2_3_1;
  wire pp_2_4_0;
  wire pp_2_4_1;
  wire pp_2_4_2;
  wire pp_2_5_0;
  wire pp_2_5_1;
  wire pp_2_6_0;
  wire pp_2_6_1;
  wire pp_2_7_0;
  wire pp_2_7_1;
  wire pp_2_8_0;
  wire pp_2_8_1;
  wire pp_2_9_0;
  wire pp_2_9_1;
  wire pp_2_9_2;
  wire pp_2_9_3;
  wire pp_2_10_0;
  wire pp_2_10_1;
  wire pp_2_10_2;
  wire pp_2_11_0;
  wire pp_2_11_1;
  wire pp_2_11_2;
  wire pp_2_12_0;
  wire pp_2_12_1;
  wire pp_2_12_2;
  wire pp_2_13_0;
  wire pp_2_13_1;
  wire pp_2_13_2;
  wire pp_2_13_3;
  wire pp_2_13_4;
  wire pp_2_14_0;
  wire pp_2_14_1;
  wire pp_2_14_2;
  wire pp_2_14_3;
  wire pp_2_15_0;
  wire pp_2_15_1;
  wire pp_2_15_2;
  wire pp_2_15_3;
  wire pp_2_16_0;
  wire pp_2_16_1;
  wire pp_2_16_2;
  wire pp_2_16_3;
  wire pp_2_17_0;
  wire pp_2_17_1;
  wire pp_2_17_2;
  wire pp_2_17_3;
  wire pp_2_18_0;
  wire pp_2_18_1;
  wire pp_2_18_2;
  wire pp_2_18_3;
  wire pp_2_18_4;
  wire pp_2_18_5;
  wire pp_2_19_0;
  wire pp_2_19_1;
  wire pp_2_19_2;
  wire pp_2_19_3;
  wire pp_2_19_4;
  wire pp_2_20_0;
  wire pp_2_20_1;
  wire pp_2_20_2;
  wire pp_2_20_3;
  wire pp_2_20_4;
  wire pp_2_21_0;
  wire pp_2_21_1;
  wire pp_2_21_2;
  wire pp_2_21_3;
  wire pp_2_21_4;
  wire pp_2_22_0;
  wire pp_2_22_1;
  wire pp_2_22_2;
  wire pp_2_22_3;
  wire pp_2_22_4;
  wire pp_2_22_5;
  wire pp_2_23_0;
  wire pp_2_23_1;
  wire pp_2_23_2;
  wire pp_2_23_3;
  wire pp_2_23_4;
  wire pp_2_23_5;
  wire pp_2_23_6;
  wire pp_2_24_0;
  wire pp_2_24_1;
  wire pp_2_24_2;
  wire pp_2_24_3;
  wire pp_2_24_4;
  wire pp_2_24_5;
  wire pp_2_24_6;
  wire pp_2_24_7;
  wire pp_2_24_8;
  wire pp_2_24_9;
  wire pp_2_24_10;
  wire pp_2_24_11;
  wire pp_2_25_0;
  wire pp_2_25_1;
  wire pp_2_25_2;
  wire pp_2_26_0;
  wire pp_2_26_1;
  wire pp_2_26_2;
  wire pp_2_26_3;
  wire pp_2_26_4;
  wire pp_2_26_5;
  wire pp_2_27_0;
  wire pp_2_27_1;
  wire pp_2_27_2;
  wire pp_2_27_3;
  wire pp_2_27_4;
  wire pp_2_27_5;
  wire pp_2_27_6;
  wire pp_2_27_7;
  wire pp_2_28_0;
  wire pp_2_28_1;
  wire pp_2_28_2;
  wire pp_2_28_3;
  wire pp_2_28_4;
  wire pp_2_28_5;
  wire pp_2_28_6;
  wire pp_2_29_0;
  wire pp_2_29_1;
  wire pp_2_29_2;
  wire pp_2_29_3;
  wire pp_2_29_4;
  wire pp_2_29_5;
  wire pp_2_29_6;
  wire pp_2_30_0;
  wire pp_2_30_1;
  wire pp_2_30_2;
  wire pp_2_30_3;
  wire pp_2_30_4;
  wire pp_2_30_5;
  wire pp_2_30_6;
  wire pp_2_31_0;
  wire pp_2_31_1;
  wire pp_2_31_2;
  wire pp_2_31_3;
  wire pp_2_31_4;
  wire pp_2_31_5;
  wire pp_2_31_6;
  wire pp_2_31_7;
  wire pp_2_32_0;
  wire pp_2_32_1;
  wire pp_2_32_2;
  wire pp_2_32_3;
  wire pp_2_32_4;
  wire pp_2_32_5;
  wire pp_2_32_6;
  wire pp_2_32_7;
  wire pp_2_32_8;
  wire pp_2_32_9;
  wire pp_2_32_10;
  wire pp_2_32_11;
  wire pp_2_33_0;
  wire pp_2_33_1;
  wire pp_2_33_2;
  wire pp_2_33_3;
  wire pp_2_33_4;
  wire pp_2_33_5;
  wire pp_2_34_0;
  wire pp_2_34_1;
  wire pp_2_34_2;
  wire pp_2_34_3;
  wire pp_2_34_4;
  wire pp_2_34_5;
  wire pp_2_34_6;
  wire pp_2_34_7;
  wire pp_2_35_0;
  wire pp_2_35_1;
  wire pp_2_35_2;
  wire pp_2_35_3;
  wire pp_2_35_4;
  wire pp_2_35_5;
  wire pp_2_35_6;
  wire pp_2_35_7;
  wire pp_2_36_0;
  wire pp_2_36_1;
  wire pp_2_36_2;
  wire pp_2_36_3;
  wire pp_2_36_4;
  wire pp_2_36_5;
  wire pp_2_36_6;
  wire pp_2_36_7;
  wire pp_2_36_8;
  wire pp_2_37_0;
  wire pp_2_37_1;
  wire pp_2_37_2;
  wire pp_2_37_3;
  wire pp_2_37_4;
  wire pp_2_37_5;
  wire pp_2_37_6;
  wire pp_2_38_0;
  wire pp_2_38_1;
  wire pp_2_38_2;
  wire pp_2_38_3;
  wire pp_2_38_4;
  wire pp_2_38_5;
  wire pp_2_38_6;
  wire pp_2_39_0;
  wire pp_2_39_1;
  wire pp_2_39_2;
  wire pp_2_39_3;
  wire pp_2_39_4;
  wire pp_2_39_5;
  wire pp_2_39_6;
  wire pp_2_39_7;
  wire pp_2_40_0;
  wire pp_2_40_1;
  wire pp_2_40_2;
  wire pp_2_40_3;
  wire pp_2_40_4;
  wire pp_2_40_5;
  wire pp_2_40_6;
  wire pp_2_40_7;
  wire pp_2_40_8;
  wire pp_2_41_0;
  wire pp_2_41_1;
  wire pp_2_41_2;
  wire pp_2_41_3;
  wire pp_2_41_4;
  wire pp_2_42_0;
  wire pp_2_42_1;
  wire pp_2_42_2;
  wire pp_2_42_3;
  wire pp_2_42_4;
  wire pp_2_42_5;
  wire pp_2_43_0;
  wire pp_2_43_1;
  wire pp_2_43_2;
  wire pp_2_43_3;
  wire pp_2_43_4;
  wire pp_2_43_5;
  wire pp_2_43_6;
  wire pp_2_44_0;
  wire pp_2_44_1;
  wire pp_2_44_2;
  wire pp_2_44_3;
  wire pp_2_44_4;
  wire pp_2_44_5;
  wire pp_2_45_0;
  wire pp_2_45_1;
  wire pp_2_45_2;
  wire pp_2_45_3;
  wire pp_2_45_4;
  wire pp_2_45_5;
  wire pp_2_45_6;
  wire pp_2_46_0;
  wire pp_2_46_1;
  wire pp_2_46_2;
  wire pp_2_46_3;
  wire pp_2_46_4;
  wire pp_2_46_5;
  wire pp_2_46_6;
  wire pp_2_47_0;
  wire pp_2_47_1;
  wire pp_2_47_2;
  wire pp_2_47_3;
  wire pp_2_47_4;
  wire pp_2_48_0;
  wire pp_2_48_1;
  wire pp_2_48_2;
  wire pp_2_48_3;
  wire pp_2_48_4;
  wire pp_2_49_0;
  wire pp_2_49_1;
  wire pp_2_49_2;
  wire pp_2_49_3;
  wire pp_2_49_4;
  wire pp_2_49_5;
  wire pp_2_50_0;
  wire pp_2_50_1;
  wire pp_2_50_2;
  wire pp_2_51_0;
  wire pp_2_51_1;
  wire pp_2_51_2;
  wire pp_2_51_3;
  wire pp_2_51_4;
  wire pp_2_52_0;
  wire pp_2_52_1;
  wire pp_2_52_2;
  wire pp_2_52_3;
  wire pp_2_53_0;
  wire pp_2_53_1;
  wire pp_2_53_2;
  wire pp_2_53_3;
  wire pp_2_53_4;
  wire pp_2_54_0;
  wire pp_2_54_1;
  wire pp_2_54_2;
  wire pp_2_54_3;
  wire pp_2_55_0;
  wire pp_2_55_1;
  wire pp_2_55_2;
  wire pp_2_55_3;
  wire pp_2_55_4;
  wire pp_2_56_0;
  wire pp_2_56_1;
  wire pp_2_56_2;
  wire pp_2_56_3;
  wire pp_2_56_4;
  wire pp_2_56_5;
  wire pp_2_57_0;
  wire pp_2_57_1;
  wire pp_2_58_0;
  wire pp_2_58_1;
  wire pp_2_58_2;
  wire pp_2_59_0;
  wire pp_2_59_1;
  wire pp_2_59_2;
  wire pp_2_59_3;
  wire pp_2_60_0;
  wire pp_2_61_0;
  wire pp_2_61_1;
  wire pp_2_61_2;
  wire pp_2_62_0;
  wire pp_2_62_1;
  wire pp_2_63_0;
  wire pp_2_63_1;
  wire pp_2_63_2;
  wire pp_3_0_0;
  wire pp_3_0_1;
  wire pp_3_1_0;
  wire pp_3_2_0;
  wire pp_3_2_1;
  wire pp_3_3_0;
  wire pp_3_3_1;
  wire pp_3_4_0;
  wire pp_3_4_1;
  wire pp_3_4_2;
  wire pp_3_5_0;
  wire pp_3_6_0;
  wire pp_3_6_1;
  wire pp_3_6_2;
  wire pp_3_7_0;
  wire pp_3_8_0;
  wire pp_3_8_1;
  wire pp_3_8_2;
  wire pp_3_9_0;
  wire pp_3_9_1;
  wire pp_3_9_2;
  wire pp_3_9_3;
  wire pp_3_10_0;
  wire pp_3_11_0;
  wire pp_3_11_1;
  wire pp_3_12_0;
  wire pp_3_12_1;
  wire pp_3_13_0;
  wire pp_3_13_1;
  wire pp_3_13_2;
  wire pp_3_13_3;
  wire pp_3_14_0;
  wire pp_3_14_1;
  wire pp_3_14_2;
  wire pp_3_15_0;
  wire pp_3_15_1;
  wire pp_3_15_2;
  wire pp_3_16_0;
  wire pp_3_16_1;
  wire pp_3_16_2;
  wire pp_3_16_3;
  wire pp_3_17_0;
  wire pp_3_17_1;
  wire pp_3_17_2;
  wire pp_3_18_0;
  wire pp_3_18_1;
  wire pp_3_18_2;
  wire pp_3_19_0;
  wire pp_3_19_1;
  wire pp_3_19_2;
  wire pp_3_19_3;
  wire pp_3_20_0;
  wire pp_3_20_1;
  wire pp_3_20_2;
  wire pp_3_20_3;
  wire pp_3_21_0;
  wire pp_3_21_1;
  wire pp_3_21_2;
  wire pp_3_21_3;
  wire pp_3_22_0;
  wire pp_3_22_1;
  wire pp_3_22_2;
  wire pp_3_22_3;
  wire pp_3_22_4;
  wire pp_3_22_5;
  wire pp_3_23_0;
  wire pp_3_23_1;
  wire pp_3_23_2;
  wire pp_3_23_3;
  wire pp_3_24_0;
  wire pp_3_24_1;
  wire pp_3_24_2;
  wire pp_3_24_3;
  wire pp_3_24_4;
  wire pp_3_24_5;
  wire pp_3_25_0;
  wire pp_3_25_1;
  wire pp_3_25_2;
  wire pp_3_25_3;
  wire pp_3_25_4;
  wire pp_3_25_5;
  wire pp_3_26_0;
  wire pp_3_26_1;
  wire pp_3_26_2;
  wire pp_3_27_0;
  wire pp_3_27_1;
  wire pp_3_27_2;
  wire pp_3_27_3;
  wire pp_3_27_4;
  wire pp_3_27_5;
  wire pp_3_28_0;
  wire pp_3_28_1;
  wire pp_3_28_2;
  wire pp_3_28_3;
  wire pp_3_28_4;
  wire pp_3_29_0;
  wire pp_3_29_1;
  wire pp_3_29_2;
  wire pp_3_29_3;
  wire pp_3_29_4;
  wire pp_3_30_0;
  wire pp_3_30_1;
  wire pp_3_30_2;
  wire pp_3_30_3;
  wire pp_3_30_4;
  wire pp_3_30_5;
  wire pp_3_31_0;
  wire pp_3_31_1;
  wire pp_3_31_2;
  wire pp_3_31_3;
  wire pp_3_31_4;
  wire pp_3_31_5;
  wire pp_3_32_0;
  wire pp_3_32_1;
  wire pp_3_32_2;
  wire pp_3_32_3;
  wire pp_3_32_4;
  wire pp_3_32_5;
  wire pp_3_33_0;
  wire pp_3_33_1;
  wire pp_3_33_2;
  wire pp_3_33_3;
  wire pp_3_33_4;
  wire pp_3_33_5;
  wire pp_3_34_0;
  wire pp_3_34_1;
  wire pp_3_34_2;
  wire pp_3_34_3;
  wire pp_3_34_4;
  wire pp_3_34_5;
  wire pp_3_35_0;
  wire pp_3_35_1;
  wire pp_3_35_2;
  wire pp_3_35_3;
  wire pp_3_35_4;
  wire pp_3_35_5;
  wire pp_3_36_0;
  wire pp_3_36_1;
  wire pp_3_36_2;
  wire pp_3_36_3;
  wire pp_3_36_4;
  wire pp_3_37_0;
  wire pp_3_37_1;
  wire pp_3_37_2;
  wire pp_3_37_3;
  wire pp_3_37_4;
  wire pp_3_37_5;
  wire pp_3_38_0;
  wire pp_3_38_1;
  wire pp_3_38_2;
  wire pp_3_38_3;
  wire pp_3_38_4;
  wire pp_3_38_5;
  wire pp_3_39_0;
  wire pp_3_39_1;
  wire pp_3_39_2;
  wire pp_3_39_3;
  wire pp_3_39_4;
  wire pp_3_39_5;
  wire pp_3_40_0;
  wire pp_3_40_1;
  wire pp_3_40_2;
  wire pp_3_40_3;
  wire pp_3_40_4;
  wire pp_3_41_0;
  wire pp_3_41_1;
  wire pp_3_41_2;
  wire pp_3_41_3;
  wire pp_3_41_4;
  wire pp_3_41_5;
  wire pp_3_42_0;
  wire pp_3_42_1;
  wire pp_3_42_2;
  wire pp_3_43_0;
  wire pp_3_43_1;
  wire pp_3_43_2;
  wire pp_3_43_3;
  wire pp_3_43_4;
  wire pp_3_44_0;
  wire pp_3_44_1;
  wire pp_3_44_2;
  wire pp_3_44_3;
  wire pp_3_44_4;
  wire pp_3_44_5;
  wire pp_3_45_0;
  wire pp_3_45_1;
  wire pp_3_45_2;
  wire pp_3_45_3;
  wire pp_3_46_0;
  wire pp_3_46_1;
  wire pp_3_46_2;
  wire pp_3_46_3;
  wire pp_3_46_4;
  wire pp_3_46_5;
  wire pp_3_46_6;
  wire pp_3_46_7;
  wire pp_3_46_8;
  wire pp_3_47_0;
  wire pp_3_47_1;
  wire pp_3_47_2;
  wire pp_3_48_0;
  wire pp_3_48_1;
  wire pp_3_48_2;
  wire pp_3_48_3;
  wire pp_3_48_4;
  wire pp_3_48_5;
  wire pp_3_49_0;
  wire pp_3_49_1;
  wire pp_3_50_0;
  wire pp_3_50_1;
  wire pp_3_50_2;
  wire pp_3_51_0;
  wire pp_3_51_1;
  wire pp_3_51_2;
  wire pp_3_51_3;
  wire pp_3_52_0;
  wire pp_3_52_1;
  wire pp_3_52_2;
  wire pp_3_53_0;
  wire pp_3_53_1;
  wire pp_3_53_2;
  wire pp_3_53_3;
  wire pp_3_54_0;
  wire pp_3_54_1;
  wire pp_3_54_2;
  wire pp_3_54_3;
  wire pp_3_54_4;
  wire pp_3_55_0;
  wire pp_3_55_1;
  wire pp_3_55_2;
  wire pp_3_56_0;
  wire pp_3_56_1;
  wire pp_3_56_2;
  wire pp_3_57_0;
  wire pp_3_57_1;
  wire pp_3_57_2;
  wire pp_3_57_3;
  wire pp_3_58_0;
  wire pp_3_58_1;
  wire pp_3_58_2;
  wire pp_3_59_0;
  wire pp_3_59_1;
  wire pp_3_59_2;
  wire pp_3_59_3;
  wire pp_3_60_0;
  wire pp_3_61_0;
  wire pp_3_62_0;
  wire pp_3_62_1;
  wire pp_3_62_2;
  wire pp_3_63_0;
  wire pp_4_0_0;
  wire pp_4_0_1;
  wire pp_4_1_0;
  wire pp_4_2_0;
  wire pp_4_2_1;
  wire pp_4_3_0;
  wire pp_4_3_1;
  wire pp_4_4_0;
  wire pp_4_4_1;
  wire pp_4_4_2;
  wire pp_4_5_0;
  wire pp_4_6_0;
  wire pp_4_6_1;
  wire pp_4_6_2;
  wire pp_4_7_0;
  wire pp_4_8_0;
  wire pp_4_8_1;
  wire pp_4_8_2;
  wire pp_4_9_0;
  wire pp_4_9_1;
  wire pp_4_10_0;
  wire pp_4_10_1;
  wire pp_4_11_0;
  wire pp_4_12_0;
  wire pp_4_12_1;
  wire pp_4_13_0;
  wire pp_4_13_1;
  wire pp_4_13_2;
  wire pp_4_14_0;
  wire pp_4_14_1;
  wire pp_4_15_0;
  wire pp_4_15_1;
  wire pp_4_16_0;
  wire pp_4_16_1;
  wire pp_4_16_2;
  wire pp_4_17_0;
  wire pp_4_17_1;
  wire pp_4_18_0;
  wire pp_4_18_1;
  wire pp_4_19_0;
  wire pp_4_19_1;
  wire pp_4_19_2;
  wire pp_4_20_0;
  wire pp_4_20_1;
  wire pp_4_20_2;
  wire pp_4_21_0;
  wire pp_4_21_1;
  wire pp_4_21_2;
  wire pp_4_22_0;
  wire pp_4_22_1;
  wire pp_4_22_2;
  wire pp_4_23_0;
  wire pp_4_23_1;
  wire pp_4_23_2;
  wire pp_4_23_3;
  wire pp_4_24_0;
  wire pp_4_24_1;
  wire pp_4_24_2;
  wire pp_4_25_0;
  wire pp_4_25_1;
  wire pp_4_25_2;
  wire pp_4_25_3;
  wire pp_4_26_0;
  wire pp_4_26_1;
  wire pp_4_26_2;
  wire pp_4_27_0;
  wire pp_4_27_1;
  wire pp_4_27_2;
  wire pp_4_28_0;
  wire pp_4_28_1;
  wire pp_4_28_2;
  wire pp_4_28_3;
  wire pp_4_28_4;
  wire pp_4_28_5;
  wire pp_4_29_0;
  wire pp_4_29_1;
  wire pp_4_29_2;
  wire pp_4_30_0;
  wire pp_4_30_1;
  wire pp_4_30_2;
  wire pp_4_30_3;
  wire pp_4_31_0;
  wire pp_4_31_1;
  wire pp_4_31_2;
  wire pp_4_31_3;
  wire pp_4_31_4;
  wire pp_4_31_5;
  wire pp_4_32_0;
  wire pp_4_32_1;
  wire pp_4_32_2;
  wire pp_4_33_0;
  wire pp_4_33_1;
  wire pp_4_33_2;
  wire pp_4_33_3;
  wire pp_4_34_0;
  wire pp_4_34_1;
  wire pp_4_34_2;
  wire pp_4_34_3;
  wire pp_4_35_0;
  wire pp_4_35_1;
  wire pp_4_35_2;
  wire pp_4_35_3;
  wire pp_4_36_0;
  wire pp_4_36_1;
  wire pp_4_36_2;
  wire pp_4_36_3;
  wire pp_4_36_4;
  wire pp_4_37_0;
  wire pp_4_37_1;
  wire pp_4_37_2;
  wire pp_4_38_0;
  wire pp_4_38_1;
  wire pp_4_38_2;
  wire pp_4_38_3;
  wire pp_4_39_0;
  wire pp_4_39_1;
  wire pp_4_39_2;
  wire pp_4_39_3;
  wire pp_4_40_0;
  wire pp_4_40_1;
  wire pp_4_40_2;
  wire pp_4_40_3;
  wire pp_4_40_4;
  wire pp_4_40_5;
  wire pp_4_41_0;
  wire pp_4_41_1;
  wire pp_4_41_2;
  wire pp_4_42_0;
  wire pp_4_42_1;
  wire pp_4_42_2;
  wire pp_4_43_0;
  wire pp_4_43_1;
  wire pp_4_43_2;
  wire pp_4_43_3;
  wire pp_4_44_0;
  wire pp_4_44_1;
  wire pp_4_44_2;
  wire pp_4_45_0;
  wire pp_4_45_1;
  wire pp_4_45_2;
  wire pp_4_45_3;
  wire pp_4_45_4;
  wire pp_4_45_5;
  wire pp_4_46_0;
  wire pp_4_46_1;
  wire pp_4_46_2;
  wire pp_4_47_0;
  wire pp_4_47_1;
  wire pp_4_47_2;
  wire pp_4_47_3;
  wire pp_4_47_4;
  wire pp_4_47_5;
  wire pp_4_48_0;
  wire pp_4_48_1;
  wire pp_4_49_0;
  wire pp_4_49_1;
  wire pp_4_49_2;
  wire pp_4_49_3;
  wire pp_4_50_0;
  wire pp_4_51_0;
  wire pp_4_51_1;
  wire pp_4_51_2;
  wire pp_4_52_0;
  wire pp_4_52_1;
  wire pp_4_53_0;
  wire pp_4_53_1;
  wire pp_4_53_2;
  wire pp_4_54_0;
  wire pp_4_54_1;
  wire pp_4_54_2;
  wire pp_4_54_3;
  wire pp_4_54_4;
  wire pp_4_54_5;
  wire pp_4_55_0;
  wire pp_4_56_0;
  wire pp_4_56_1;
  wire pp_4_57_0;
  wire pp_4_57_1;
  wire pp_4_57_2;
  wire pp_4_58_0;
  wire pp_4_58_1;
  wire pp_4_59_0;
  wire pp_4_59_1;
  wire pp_4_59_2;
  wire pp_4_60_0;
  wire pp_4_60_1;
  wire pp_4_61_0;
  wire pp_4_62_0;
  wire pp_4_62_1;
  wire pp_4_62_2;
  wire pp_4_63_0;
  wire pp_5_0_0;
  wire pp_5_0_1;
  wire pp_5_1_0;
  wire pp_5_2_0;
  wire pp_5_2_1;
  wire pp_5_3_0;
  wire pp_5_3_1;
  wire pp_5_4_0;
  wire pp_5_4_1;
  wire pp_5_5_0;
  wire pp_5_5_1;
  wire pp_5_6_0;
  wire pp_5_6_1;
  wire pp_5_7_0;
  wire pp_5_7_1;
  wire pp_5_8_0;
  wire pp_5_8_1;
  wire pp_5_8_2;
  wire pp_5_9_0;
  wire pp_5_10_0;
  wire pp_5_10_1;
  wire pp_5_11_0;
  wire pp_5_11_1;
  wire pp_5_12_0;
  wire pp_5_12_1;
  wire pp_5_13_0;
  wire pp_5_13_1;
  wire pp_5_13_2;
  wire pp_5_14_0;
  wire pp_5_15_0;
  wire pp_5_15_1;
  wire pp_5_15_2;
  wire pp_5_16_0;
  wire pp_5_17_0;
  wire pp_5_17_1;
  wire pp_5_17_2;
  wire pp_5_18_0;
  wire pp_5_19_0;
  wire pp_5_19_1;
  wire pp_5_19_2;
  wire pp_5_19_3;
  wire pp_5_20_0;
  wire pp_5_21_0;
  wire pp_5_21_1;
  wire pp_5_21_2;
  wire pp_5_21_3;
  wire pp_5_22_0;
  wire pp_5_23_0;
  wire pp_5_23_1;
  wire pp_5_23_2;
  wire pp_5_23_3;
  wire pp_5_24_0;
  wire pp_5_24_1;
  wire pp_5_24_2;
  wire pp_5_25_0;
  wire pp_5_25_1;
  wire pp_5_25_2;
  wire pp_5_26_0;
  wire pp_5_26_1;
  wire pp_5_27_0;
  wire pp_5_27_1;
  wire pp_5_28_0;
  wire pp_5_28_1;
  wire pp_5_28_2;
  wire pp_5_29_0;
  wire pp_5_29_1;
  wire pp_5_29_2;
  wire pp_5_30_0;
  wire pp_5_30_1;
  wire pp_5_30_2;
  wire pp_5_31_0;
  wire pp_5_31_1;
  wire pp_5_31_2;
  wire pp_5_32_0;
  wire pp_5_32_1;
  wire pp_5_32_2;
  wire pp_5_33_0;
  wire pp_5_33_1;
  wire pp_5_33_2;
  wire pp_5_34_0;
  wire pp_5_34_1;
  wire pp_5_34_2;
  wire pp_5_35_0;
  wire pp_5_35_1;
  wire pp_5_35_2;
  wire pp_5_36_0;
  wire pp_5_36_1;
  wire pp_5_36_2;
  wire pp_5_37_0;
  wire pp_5_37_1;
  wire pp_5_37_2;
  wire pp_5_38_0;
  wire pp_5_38_1;
  wire pp_5_38_2;
  wire pp_5_39_0;
  wire pp_5_39_1;
  wire pp_5_39_2;
  wire pp_5_40_0;
  wire pp_5_40_1;
  wire pp_5_40_2;
  wire pp_5_41_0;
  wire pp_5_41_1;
  wire pp_5_41_2;
  wire pp_5_42_0;
  wire pp_5_42_1;
  wire pp_5_42_2;
  wire pp_5_43_0;
  wire pp_5_43_1;
  wire pp_5_43_2;
  wire pp_5_44_0;
  wire pp_5_44_1;
  wire pp_5_45_0;
  wire pp_5_45_1;
  wire pp_5_45_2;
  wire pp_5_46_0;
  wire pp_5_46_1;
  wire pp_5_46_2;
  wire pp_5_47_0;
  wire pp_5_47_1;
  wire pp_5_47_2;
  wire pp_5_48_0;
  wire pp_5_48_1;
  wire pp_5_48_2;
  wire pp_5_49_0;
  wire pp_5_49_1;
  wire pp_5_49_2;
  wire pp_5_50_0;
  wire pp_5_50_1;
  wire pp_5_51_0;
  wire pp_5_51_1;
  wire pp_5_51_2;
  wire pp_5_52_0;
  wire pp_5_53_0;
  wire pp_5_53_1;
  wire pp_5_53_2;
  wire pp_5_53_3;
  wire pp_5_54_0;
  wire pp_5_54_1;
  wire pp_5_55_0;
  wire pp_5_55_1;
  wire pp_5_55_2;
  wire pp_5_56_0;
  wire pp_5_56_1;
  wire pp_5_57_0;
  wire pp_5_57_1;
  wire pp_5_57_2;
  wire pp_5_58_0;
  wire pp_5_58_1;
  wire pp_5_59_0;
  wire pp_5_60_0;
  wire pp_5_60_1;
  wire pp_5_60_2;
  wire pp_5_61_0;
  wire pp_5_62_0;
  wire pp_5_62_1;
  wire pp_5_62_2;
  wire pp_5_63_0;
  wire pp_6_0_0;
  wire pp_6_0_1;
  wire pp_6_1_0;
  wire pp_6_2_0;
  wire pp_6_2_1;
  wire pp_6_3_0;
  wire pp_6_3_1;
  wire pp_6_4_0;
  wire pp_6_4_1;
  wire pp_6_5_0;
  wire pp_6_5_1;
  wire pp_6_6_0;
  wire pp_6_6_1;
  wire pp_6_7_0;
  wire pp_6_7_1;
  wire pp_6_8_0;
  wire pp_6_8_1;
  wire pp_6_9_0;
  wire pp_6_9_1;
  wire pp_6_10_0;
  wire pp_6_10_1;
  wire pp_6_11_0;
  wire pp_6_11_1;
  wire pp_6_12_0;
  wire pp_6_12_1;
  wire pp_6_13_0;
  wire pp_6_13_1;
  wire pp_6_14_0;
  wire pp_6_14_1;
  wire pp_6_15_0;
  wire pp_6_15_1;
  wire pp_6_16_0;
  wire pp_6_16_1;
  wire pp_6_17_0;
  wire pp_6_17_1;
  wire pp_6_18_0;
  wire pp_6_18_1;
  wire pp_6_19_0;
  wire pp_6_19_1;
  wire pp_6_20_0;
  wire pp_6_20_1;
  wire pp_6_21_0;
  wire pp_6_21_1;
  wire pp_6_22_0;
  wire pp_6_22_1;
  wire pp_6_23_0;
  wire pp_6_23_1;
  wire pp_6_24_0;
  wire pp_6_24_1;
  wire pp_6_25_0;
  wire pp_6_25_1;
  wire pp_6_26_0;
  wire pp_6_26_1;
  wire pp_6_27_0;
  wire pp_6_27_1;
  wire pp_6_28_0;
  wire pp_6_28_1;
  wire pp_6_29_0;
  wire pp_6_29_1;
  wire pp_6_30_0;
  wire pp_6_30_1;
  wire pp_6_31_0;
  wire pp_6_31_1;
  wire pp_6_32_0;
  wire pp_6_32_1;
  wire pp_6_33_0;
  wire pp_6_33_1;
  wire pp_6_34_0;
  wire pp_6_34_1;
  wire pp_6_35_0;
  wire pp_6_35_1;
  wire pp_6_36_0;
  wire pp_6_36_1;
  wire pp_6_37_0;
  wire pp_6_37_1;
  wire pp_6_38_0;
  wire pp_6_38_1;
  wire pp_6_39_0;
  wire pp_6_39_1;
  wire pp_6_40_0;
  wire pp_6_40_1;
  wire pp_6_41_0;
  wire pp_6_41_1;
  wire pp_6_42_0;
  wire pp_6_42_1;
  wire pp_6_43_0;
  wire pp_6_43_1;
  wire pp_6_44_0;
  wire pp_6_44_1;
  wire pp_6_45_0;
  wire pp_6_45_1;
  wire pp_6_46_0;
  wire pp_6_46_1;
  wire pp_6_47_0;
  wire pp_6_47_1;
  wire pp_6_48_0;
  wire pp_6_48_1;
  wire pp_6_49_0;
  wire pp_6_49_1;
  wire pp_6_50_0;
  wire pp_6_50_1;
  wire pp_6_51_0;
  wire pp_6_51_1;
  wire pp_6_52_0;
  wire pp_6_52_1;
  wire pp_6_53_0;
  wire pp_6_53_1;
  wire pp_6_54_0;
  wire pp_6_54_1;
  wire pp_6_55_0;
  wire pp_6_55_1;
  wire pp_6_56_0;
  wire pp_6_56_1;
  wire pp_6_57_0;
  wire pp_6_57_1;
  wire pp_6_58_0;
  wire pp_6_58_1;
  wire pp_6_59_0;
  wire pp_6_59_1;
  wire pp_6_60_0;
  wire pp_6_60_1;
  wire pp_6_61_0;
  wire pp_6_61_1;
  wire pp_6_62_0;
  wire pp_6_62_1;
  wire pp_6_63_0;
  wire pp_6_63_1;
  assign pp_0_0_0 = pp_0_0;
  assign pp_0_0_1 = be_c_0;
  assign pp_0_1_0 = pp_0_1;
  assign pp_0_2_0 = pp_0_2;
  assign pp_0_2_1 = pp_1_2;
  assign pp_0_2_2 = be_c_1;
  assign pp_0_3_0 = pp_0_3;
  assign pp_0_3_1 = pp_1_3;
  assign pp_0_4_0 = pp_0_4;
  assign pp_0_4_1 = pp_1_4;
  assign pp_0_4_2 = pp_2_4;
  assign pp_0_4_3 = be_c_2;
  assign pp_0_5_0 = pp_0_5;
  assign pp_0_5_1 = pp_1_5;
  assign pp_0_5_2 = pp_2_5;
  assign pp_0_6_0 = pp_0_6;
  assign pp_0_6_1 = pp_1_6;
  assign pp_0_6_2 = pp_2_6;
  assign pp_0_6_3 = pp_3_6;
  assign pp_0_6_4 = be_c_3;
  assign pp_0_7_0 = pp_0_7;
  assign pp_0_7_1 = pp_1_7;
  assign pp_0_7_2 = pp_2_7;
  assign pp_0_7_3 = pp_3_7;
  assign pp_0_8_0 = pp_0_8;
  assign pp_0_8_1 = pp_1_8;
  assign pp_0_8_2 = pp_2_8;
  assign pp_0_8_3 = pp_3_8;
  assign pp_0_8_4 = pp_4_8;
  assign pp_0_8_5 = be_c_4;
  assign pp_0_9_0 = pp_0_9;
  assign pp_0_9_1 = pp_1_9;
  assign pp_0_9_2 = pp_2_9;
  assign pp_0_9_3 = pp_3_9;
  assign pp_0_9_4 = pp_4_9;
  assign pp_0_10_0 = pp_0_10;
  assign pp_0_10_1 = pp_1_10;
  assign pp_0_10_2 = pp_2_10;
  assign pp_0_10_3 = pp_3_10;
  assign pp_0_10_4 = pp_4_10;
  assign pp_0_10_5 = pp_5_10;
  assign pp_0_10_6 = be_c_5;
  assign pp_0_11_0 = pp_0_11;
  assign pp_0_11_1 = pp_1_11;
  assign pp_0_11_2 = pp_2_11;
  assign pp_0_11_3 = pp_3_11;
  assign pp_0_11_4 = pp_4_11;
  assign pp_0_11_5 = pp_5_11;
  assign pp_0_12_0 = pp_0_12;
  assign pp_0_12_1 = pp_1_12;
  assign pp_0_12_2 = pp_2_12;
  assign pp_0_12_3 = pp_3_12;
  assign pp_0_12_4 = pp_4_12;
  assign pp_0_12_5 = pp_5_12;
  assign pp_0_12_6 = pp_6_12;
  assign pp_0_12_7 = be_c_6;
  assign pp_0_13_0 = pp_0_13;
  assign pp_0_13_1 = pp_1_13;
  assign pp_0_13_2 = pp_2_13;
  assign pp_0_13_3 = pp_3_13;
  assign pp_0_13_4 = pp_4_13;
  assign pp_0_13_5 = pp_5_13;
  assign pp_0_13_6 = pp_6_13;
  assign pp_0_14_0 = pp_0_14;
  assign pp_0_14_1 = pp_1_14;
  assign pp_0_14_2 = pp_2_14;
  assign pp_0_14_3 = pp_3_14;
  assign pp_0_14_4 = pp_4_14;
  assign pp_0_14_5 = pp_5_14;
  assign pp_0_14_6 = pp_6_14;
  assign pp_0_14_7 = pp_7_14;
  assign pp_0_14_8 = be_c_7;
  assign pp_0_15_0 = pp_0_15;
  assign pp_0_15_1 = pp_1_15;
  assign pp_0_15_2 = pp_2_15;
  assign pp_0_15_3 = pp_3_15;
  assign pp_0_15_4 = pp_4_15;
  assign pp_0_15_5 = pp_5_15;
  assign pp_0_15_6 = pp_6_15;
  assign pp_0_15_7 = pp_7_15;
  assign pp_0_16_0 = pp_0_16;
  assign pp_0_16_1 = pp_1_16;
  assign pp_0_16_2 = pp_2_16;
  assign pp_0_16_3 = pp_3_16;
  assign pp_0_16_4 = pp_4_16;
  assign pp_0_16_5 = pp_5_16;
  assign pp_0_16_6 = pp_6_16;
  assign pp_0_16_7 = pp_7_16;
  assign pp_0_16_8 = pp_8_16;
  assign pp_0_16_9 = be_c_8;
  assign pp_0_17_0 = pp_0_17;
  assign pp_0_17_1 = pp_1_17;
  assign pp_0_17_2 = pp_2_17;
  assign pp_0_17_3 = pp_3_17;
  assign pp_0_17_4 = pp_4_17;
  assign pp_0_17_5 = pp_5_17;
  assign pp_0_17_6 = pp_6_17;
  assign pp_0_17_7 = pp_7_17;
  assign pp_0_17_8 = pp_8_17;
  assign pp_0_18_0 = pp_0_18;
  assign pp_0_18_1 = pp_1_18;
  assign pp_0_18_2 = pp_2_18;
  assign pp_0_18_3 = pp_3_18;
  assign pp_0_18_4 = pp_4_18;
  assign pp_0_18_5 = pp_5_18;
  assign pp_0_18_6 = pp_6_18;
  assign pp_0_18_7 = pp_7_18;
  assign pp_0_18_8 = pp_8_18;
  assign pp_0_18_9 = pp_9_18;
  assign pp_0_18_10 = be_c_9;
  assign pp_0_19_0 = pp_0_19;
  assign pp_0_19_1 = pp_1_19;
  assign pp_0_19_2 = pp_2_19;
  assign pp_0_19_3 = pp_3_19;
  assign pp_0_19_4 = pp_4_19;
  assign pp_0_19_5 = pp_5_19;
  assign pp_0_19_6 = pp_6_19;
  assign pp_0_19_7 = pp_7_19;
  assign pp_0_19_8 = pp_8_19;
  assign pp_0_19_9 = pp_9_19;
  assign pp_0_20_0 = pp_0_20;
  assign pp_0_20_1 = pp_1_20;
  assign pp_0_20_2 = pp_2_20;
  assign pp_0_20_3 = pp_3_20;
  assign pp_0_20_4 = pp_4_20;
  assign pp_0_20_5 = pp_5_20;
  assign pp_0_20_6 = pp_6_20;
  assign pp_0_20_7 = pp_7_20;
  assign pp_0_20_8 = pp_8_20;
  assign pp_0_20_9 = pp_9_20;
  assign pp_0_20_10 = pp_10_20;
  assign pp_0_20_11 = be_c_10;
  assign pp_0_21_0 = pp_0_21;
  assign pp_0_21_1 = pp_1_21;
  assign pp_0_21_2 = pp_2_21;
  assign pp_0_21_3 = pp_3_21;
  assign pp_0_21_4 = pp_4_21;
  assign pp_0_21_5 = pp_5_21;
  assign pp_0_21_6 = pp_6_21;
  assign pp_0_21_7 = pp_7_21;
  assign pp_0_21_8 = pp_8_21;
  assign pp_0_21_9 = pp_9_21;
  assign pp_0_21_10 = pp_10_21;
  assign pp_0_22_0 = pp_0_22;
  assign pp_0_22_1 = pp_1_22;
  assign pp_0_22_2 = pp_2_22;
  assign pp_0_22_3 = pp_3_22;
  assign pp_0_22_4 = pp_4_22;
  assign pp_0_22_5 = pp_5_22;
  assign pp_0_22_6 = pp_6_22;
  assign pp_0_22_7 = pp_7_22;
  assign pp_0_22_8 = pp_8_22;
  assign pp_0_22_9 = pp_9_22;
  assign pp_0_22_10 = pp_10_22;
  assign pp_0_22_11 = pp_11_22;
  assign pp_0_22_12 = be_c_11;
  assign pp_0_23_0 = pp_0_23;
  assign pp_0_23_1 = pp_1_23;
  assign pp_0_23_2 = pp_2_23;
  assign pp_0_23_3 = pp_3_23;
  assign pp_0_23_4 = pp_4_23;
  assign pp_0_23_5 = pp_5_23;
  assign pp_0_23_6 = pp_6_23;
  assign pp_0_23_7 = pp_7_23;
  assign pp_0_23_8 = pp_8_23;
  assign pp_0_23_9 = pp_9_23;
  assign pp_0_23_10 = pp_10_23;
  assign pp_0_23_11 = pp_11_23;
  assign pp_0_24_0 = pp_0_24;
  assign pp_0_24_1 = pp_1_24;
  assign pp_0_24_2 = pp_2_24;
  assign pp_0_24_3 = pp_3_24;
  assign pp_0_24_4 = pp_4_24;
  assign pp_0_24_5 = pp_5_24;
  assign pp_0_24_6 = pp_6_24;
  assign pp_0_24_7 = pp_7_24;
  assign pp_0_24_8 = pp_8_24;
  assign pp_0_24_9 = pp_9_24;
  assign pp_0_24_10 = pp_10_24;
  assign pp_0_24_11 = pp_11_24;
  assign pp_0_24_12 = pp_12_24;
  assign pp_0_24_13 = be_c_12;
  assign pp_0_25_0 = pp_0_25;
  assign pp_0_25_1 = pp_1_25;
  assign pp_0_25_2 = pp_2_25;
  assign pp_0_25_3 = pp_3_25;
  assign pp_0_25_4 = pp_4_25;
  assign pp_0_25_5 = pp_5_25;
  assign pp_0_25_6 = pp_6_25;
  assign pp_0_25_7 = pp_7_25;
  assign pp_0_25_8 = pp_8_25;
  assign pp_0_25_9 = pp_9_25;
  assign pp_0_25_10 = pp_10_25;
  assign pp_0_25_11 = pp_11_25;
  assign pp_0_25_12 = pp_12_25;
  assign pp_0_26_0 = pp_0_26;
  assign pp_0_26_1 = pp_1_26;
  assign pp_0_26_2 = pp_2_26;
  assign pp_0_26_3 = pp_3_26;
  assign pp_0_26_4 = pp_4_26;
  assign pp_0_26_5 = pp_5_26;
  assign pp_0_26_6 = pp_6_26;
  assign pp_0_26_7 = pp_7_26;
  assign pp_0_26_8 = pp_8_26;
  assign pp_0_26_9 = pp_9_26;
  assign pp_0_26_10 = pp_10_26;
  assign pp_0_26_11 = pp_11_26;
  assign pp_0_26_12 = pp_12_26;
  assign pp_0_26_13 = pp_13_26;
  assign pp_0_26_14 = be_c_13;
  assign pp_0_27_0 = pp_0_27;
  assign pp_0_27_1 = pp_1_27;
  assign pp_0_27_2 = pp_2_27;
  assign pp_0_27_3 = pp_3_27;
  assign pp_0_27_4 = pp_4_27;
  assign pp_0_27_5 = pp_5_27;
  assign pp_0_27_6 = pp_6_27;
  assign pp_0_27_7 = pp_7_27;
  assign pp_0_27_8 = pp_8_27;
  assign pp_0_27_9 = pp_9_27;
  assign pp_0_27_10 = pp_10_27;
  assign pp_0_27_11 = pp_11_27;
  assign pp_0_27_12 = pp_12_27;
  assign pp_0_27_13 = pp_13_27;
  assign pp_0_28_0 = pp_0_28;
  assign pp_0_28_1 = pp_1_28;
  assign pp_0_28_2 = pp_2_28;
  assign pp_0_28_3 = pp_3_28;
  assign pp_0_28_4 = pp_4_28;
  assign pp_0_28_5 = pp_5_28;
  assign pp_0_28_6 = pp_6_28;
  assign pp_0_28_7 = pp_7_28;
  assign pp_0_28_8 = pp_8_28;
  assign pp_0_28_9 = pp_9_28;
  assign pp_0_28_10 = pp_10_28;
  assign pp_0_28_11 = pp_11_28;
  assign pp_0_28_12 = pp_12_28;
  assign pp_0_28_13 = pp_13_28;
  assign pp_0_28_14 = pp_14_28;
  assign pp_0_28_15 = be_c_14;
  assign pp_0_29_0 = pp_0_29;
  assign pp_0_29_1 = pp_1_29;
  assign pp_0_29_2 = pp_2_29;
  assign pp_0_29_3 = pp_3_29;
  assign pp_0_29_4 = pp_4_29;
  assign pp_0_29_5 = pp_5_29;
  assign pp_0_29_6 = pp_6_29;
  assign pp_0_29_7 = pp_7_29;
  assign pp_0_29_8 = pp_8_29;
  assign pp_0_29_9 = pp_9_29;
  assign pp_0_29_10 = pp_10_29;
  assign pp_0_29_11 = pp_11_29;
  assign pp_0_29_12 = pp_12_29;
  assign pp_0_29_13 = pp_13_29;
  assign pp_0_29_14 = pp_14_29;
  assign pp_0_30_0 = pp_0_30;
  assign pp_0_30_1 = pp_1_30;
  assign pp_0_30_2 = pp_2_30;
  assign pp_0_30_3 = pp_3_30;
  assign pp_0_30_4 = pp_4_30;
  assign pp_0_30_5 = pp_5_30;
  assign pp_0_30_6 = pp_6_30;
  assign pp_0_30_7 = pp_7_30;
  assign pp_0_30_8 = pp_8_30;
  assign pp_0_30_9 = pp_9_30;
  assign pp_0_30_10 = pp_10_30;
  assign pp_0_30_11 = pp_11_30;
  assign pp_0_30_12 = pp_12_30;
  assign pp_0_30_13 = pp_13_30;
  assign pp_0_30_14 = pp_14_30;
  assign pp_0_30_15 = pp_15_30;
  assign pp_0_30_16 = be_c_15;
  assign pp_0_31_0 = pp_0_31;
  assign pp_0_31_1 = pp_1_31;
  assign pp_0_31_2 = pp_2_31;
  assign pp_0_31_3 = pp_3_31;
  assign pp_0_31_4 = pp_4_31;
  assign pp_0_31_5 = pp_5_31;
  assign pp_0_31_6 = pp_6_31;
  assign pp_0_31_7 = pp_7_31;
  assign pp_0_31_8 = pp_8_31;
  assign pp_0_31_9 = pp_9_31;
  assign pp_0_31_10 = pp_10_31;
  assign pp_0_31_11 = pp_11_31;
  assign pp_0_31_12 = pp_12_31;
  assign pp_0_31_13 = pp_13_31;
  assign pp_0_31_14 = pp_14_31;
  assign pp_0_31_15 = pp_15_31;
  assign pp_0_32_0 = pp_0_32;
  assign pp_0_32_1 = pp_1_32;
  assign pp_0_32_2 = pp_2_32;
  assign pp_0_32_3 = pp_3_32;
  assign pp_0_32_4 = pp_4_32;
  assign pp_0_32_5 = pp_5_32;
  assign pp_0_32_6 = pp_6_32;
  assign pp_0_32_7 = pp_7_32;
  assign pp_0_32_8 = pp_8_32;
  assign pp_0_32_9 = pp_9_32;
  assign pp_0_32_10 = pp_10_32;
  assign pp_0_32_11 = pp_11_32;
  assign pp_0_32_12 = pp_12_32;
  assign pp_0_32_13 = pp_13_32;
  assign pp_0_32_14 = pp_14_32;
  assign pp_0_32_15 = pp_15_32;
  assign pp_0_32_16 = pp_16_32;
  assign pp_0_33_0 = pp_0_33;
  assign pp_0_33_1 = pp_1_33;
  assign pp_0_33_2 = pp_2_33;
  assign pp_0_33_3 = pp_3_33;
  assign pp_0_33_4 = pp_4_33;
  assign pp_0_33_5 = pp_5_33;
  assign pp_0_33_6 = pp_6_33;
  assign pp_0_33_7 = pp_7_33;
  assign pp_0_33_8 = pp_8_33;
  assign pp_0_33_9 = pp_9_33;
  assign pp_0_33_10 = pp_10_33;
  assign pp_0_33_11 = pp_11_33;
  assign pp_0_33_12 = pp_12_33;
  assign pp_0_33_13 = pp_13_33;
  assign pp_0_33_14 = pp_14_33;
  assign pp_0_33_15 = pp_15_33;
  assign pp_0_33_16 = pp_16_33;
  assign pp_0_34_0 = pp_0_33;
  assign pp_0_34_1 = pp_1_34;
  assign pp_0_34_2 = pp_2_34;
  assign pp_0_34_3 = pp_3_34;
  assign pp_0_34_4 = pp_4_34;
  assign pp_0_34_5 = pp_5_34;
  assign pp_0_34_6 = pp_6_34;
  assign pp_0_34_7 = pp_7_34;
  assign pp_0_34_8 = pp_8_34;
  assign pp_0_34_9 = pp_9_34;
  assign pp_0_34_10 = pp_10_34;
  assign pp_0_34_11 = pp_11_34;
  assign pp_0_34_12 = pp_12_34;
  assign pp_0_34_13 = pp_13_34;
  assign pp_0_34_14 = pp_14_34;
  assign pp_0_34_15 = pp_15_34;
  assign pp_0_34_16 = pp_16_34;
  assign pp_0_35_0 = not_pp_0_35;
  assign pp_0_35_1 = not_pp_1_35;
  assign pp_0_35_2 = pp_2_35;
  assign pp_0_35_3 = pp_3_35;
  assign pp_0_35_4 = pp_4_35;
  assign pp_0_35_5 = pp_5_35;
  assign pp_0_35_6 = pp_6_35;
  assign pp_0_35_7 = pp_7_35;
  assign pp_0_35_8 = pp_8_35;
  assign pp_0_35_9 = pp_9_35;
  assign pp_0_35_10 = pp_10_35;
  assign pp_0_35_11 = pp_11_35;
  assign pp_0_35_12 = pp_12_35;
  assign pp_0_35_13 = pp_13_35;
  assign pp_0_35_14 = pp_14_35;
  assign pp_0_35_15 = pp_15_35;
  assign pp_0_35_16 = pp_16_35;
  assign pp_0_36_0 = one;
  assign pp_0_36_1 = pp_2_36;
  assign pp_0_36_2 = pp_3_36;
  assign pp_0_36_3 = pp_4_36;
  assign pp_0_36_4 = pp_5_36;
  assign pp_0_36_5 = pp_6_36;
  assign pp_0_36_6 = pp_7_36;
  assign pp_0_36_7 = pp_8_36;
  assign pp_0_36_8 = pp_9_36;
  assign pp_0_36_9 = pp_10_36;
  assign pp_0_36_10 = pp_11_36;
  assign pp_0_36_11 = pp_12_36;
  assign pp_0_36_12 = pp_13_36;
  assign pp_0_36_13 = pp_14_36;
  assign pp_0_36_14 = pp_15_36;
  assign pp_0_36_15 = pp_16_36;
  assign pp_0_37_0 = not_pp_2_37;
  assign pp_0_37_1 = pp_3_37;
  assign pp_0_37_2 = pp_4_37;
  assign pp_0_37_3 = pp_5_37;
  assign pp_0_37_4 = pp_6_37;
  assign pp_0_37_5 = pp_7_37;
  assign pp_0_37_6 = pp_8_37;
  assign pp_0_37_7 = pp_9_37;
  assign pp_0_37_8 = pp_10_37;
  assign pp_0_37_9 = pp_11_37;
  assign pp_0_37_10 = pp_12_37;
  assign pp_0_37_11 = pp_13_37;
  assign pp_0_37_12 = pp_14_37;
  assign pp_0_37_13 = pp_15_37;
  assign pp_0_37_14 = pp_16_37;
  assign pp_0_38_0 = one;
  assign pp_0_38_1 = pp_3_38;
  assign pp_0_38_2 = pp_4_38;
  assign pp_0_38_3 = pp_5_38;
  assign pp_0_38_4 = pp_6_38;
  assign pp_0_38_5 = pp_7_38;
  assign pp_0_38_6 = pp_8_38;
  assign pp_0_38_7 = pp_9_38;
  assign pp_0_38_8 = pp_10_38;
  assign pp_0_38_9 = pp_11_38;
  assign pp_0_38_10 = pp_12_38;
  assign pp_0_38_11 = pp_13_38;
  assign pp_0_38_12 = pp_14_38;
  assign pp_0_38_13 = pp_15_38;
  assign pp_0_38_14 = pp_16_38;
  assign pp_0_39_0 = not_pp_3_39;
  assign pp_0_39_1 = pp_4_39;
  assign pp_0_39_2 = pp_5_39;
  assign pp_0_39_3 = pp_6_39;
  assign pp_0_39_4 = pp_7_39;
  assign pp_0_39_5 = pp_8_39;
  assign pp_0_39_6 = pp_9_39;
  assign pp_0_39_7 = pp_10_39;
  assign pp_0_39_8 = pp_11_39;
  assign pp_0_39_9 = pp_12_39;
  assign pp_0_39_10 = pp_13_39;
  assign pp_0_39_11 = pp_14_39;
  assign pp_0_39_12 = pp_15_39;
  assign pp_0_39_13 = pp_16_39;
  assign pp_0_40_0 = one;
  assign pp_0_40_1 = pp_4_40;
  assign pp_0_40_2 = pp_5_40;
  assign pp_0_40_3 = pp_6_40;
  assign pp_0_40_4 = pp_7_40;
  assign pp_0_40_5 = pp_8_40;
  assign pp_0_40_6 = pp_9_40;
  assign pp_0_40_7 = pp_10_40;
  assign pp_0_40_8 = pp_11_40;
  assign pp_0_40_9 = pp_12_40;
  assign pp_0_40_10 = pp_13_40;
  assign pp_0_40_11 = pp_14_40;
  assign pp_0_40_12 = pp_15_40;
  assign pp_0_40_13 = pp_16_40;
  assign pp_0_41_0 = not_pp_4_41;
  assign pp_0_41_1 = pp_5_41;
  assign pp_0_41_2 = pp_6_41;
  assign pp_0_41_3 = pp_7_41;
  assign pp_0_41_4 = pp_8_41;
  assign pp_0_41_5 = pp_9_41;
  assign pp_0_41_6 = pp_10_41;
  assign pp_0_41_7 = pp_11_41;
  assign pp_0_41_8 = pp_12_41;
  assign pp_0_41_9 = pp_13_41;
  assign pp_0_41_10 = pp_14_41;
  assign pp_0_41_11 = pp_15_41;
  assign pp_0_41_12 = pp_16_41;
  assign pp_0_42_0 = one;
  assign pp_0_42_1 = pp_5_42;
  assign pp_0_42_2 = pp_6_42;
  assign pp_0_42_3 = pp_7_42;
  assign pp_0_42_4 = pp_8_42;
  assign pp_0_42_5 = pp_9_42;
  assign pp_0_42_6 = pp_10_42;
  assign pp_0_42_7 = pp_11_42;
  assign pp_0_42_8 = pp_12_42;
  assign pp_0_42_9 = pp_13_42;
  assign pp_0_42_10 = pp_14_42;
  assign pp_0_42_11 = pp_15_42;
  assign pp_0_42_12 = pp_16_42;
  assign pp_0_43_0 = not_pp_5_43;
  assign pp_0_43_1 = pp_6_43;
  assign pp_0_43_2 = pp_7_43;
  assign pp_0_43_3 = pp_8_43;
  assign pp_0_43_4 = pp_9_43;
  assign pp_0_43_5 = pp_10_43;
  assign pp_0_43_6 = pp_11_43;
  assign pp_0_43_7 = pp_12_43;
  assign pp_0_43_8 = pp_13_43;
  assign pp_0_43_9 = pp_14_43;
  assign pp_0_43_10 = pp_15_43;
  assign pp_0_43_11 = pp_16_43;
  assign pp_0_44_0 = one;
  assign pp_0_44_1 = pp_6_44;
  assign pp_0_44_2 = pp_7_44;
  assign pp_0_44_3 = pp_8_44;
  assign pp_0_44_4 = pp_9_44;
  assign pp_0_44_5 = pp_10_44;
  assign pp_0_44_6 = pp_11_44;
  assign pp_0_44_7 = pp_12_44;
  assign pp_0_44_8 = pp_13_44;
  assign pp_0_44_9 = pp_14_44;
  assign pp_0_44_10 = pp_15_44;
  assign pp_0_44_11 = pp_16_44;
  assign pp_0_45_0 = not_pp_6_45;
  assign pp_0_45_1 = pp_7_45;
  assign pp_0_45_2 = pp_8_45;
  assign pp_0_45_3 = pp_9_45;
  assign pp_0_45_4 = pp_10_45;
  assign pp_0_45_5 = pp_11_45;
  assign pp_0_45_6 = pp_12_45;
  assign pp_0_45_7 = pp_13_45;
  assign pp_0_45_8 = pp_14_45;
  assign pp_0_45_9 = pp_15_45;
  assign pp_0_45_10 = pp_16_45;
  assign pp_0_46_0 = one;
  assign pp_0_46_1 = pp_7_46;
  assign pp_0_46_2 = pp_8_46;
  assign pp_0_46_3 = pp_9_46;
  assign pp_0_46_4 = pp_10_46;
  assign pp_0_46_5 = pp_11_46;
  assign pp_0_46_6 = pp_12_46;
  assign pp_0_46_7 = pp_13_46;
  assign pp_0_46_8 = pp_14_46;
  assign pp_0_46_9 = pp_15_46;
  assign pp_0_46_10 = pp_16_46;
  assign pp_0_47_0 = not_pp_7_47;
  assign pp_0_47_1 = pp_8_47;
  assign pp_0_47_2 = pp_9_47;
  assign pp_0_47_3 = pp_10_47;
  assign pp_0_47_4 = pp_11_47;
  assign pp_0_47_5 = pp_12_47;
  assign pp_0_47_6 = pp_13_47;
  assign pp_0_47_7 = pp_14_47;
  assign pp_0_47_8 = pp_15_47;
  assign pp_0_47_9 = pp_16_47;
  assign pp_0_48_0 = one;
  assign pp_0_48_1 = pp_8_48;
  assign pp_0_48_2 = pp_9_48;
  assign pp_0_48_3 = pp_10_48;
  assign pp_0_48_4 = pp_11_48;
  assign pp_0_48_5 = pp_12_48;
  assign pp_0_48_6 = pp_13_48;
  assign pp_0_48_7 = pp_14_48;
  assign pp_0_48_8 = pp_15_48;
  assign pp_0_48_9 = pp_16_48;
  assign pp_0_49_0 = not_pp_8_49;
  assign pp_0_49_1 = pp_9_49;
  assign pp_0_49_2 = pp_10_49;
  assign pp_0_49_3 = pp_11_49;
  assign pp_0_49_4 = pp_12_49;
  assign pp_0_49_5 = pp_13_49;
  assign pp_0_49_6 = pp_14_49;
  assign pp_0_49_7 = pp_15_49;
  assign pp_0_49_8 = pp_16_49;
  assign pp_0_50_0 = one;
  assign pp_0_50_1 = pp_9_50;
  assign pp_0_50_2 = pp_10_50;
  assign pp_0_50_3 = pp_11_50;
  assign pp_0_50_4 = pp_12_50;
  assign pp_0_50_5 = pp_13_50;
  assign pp_0_50_6 = pp_14_50;
  assign pp_0_50_7 = pp_15_50;
  assign pp_0_50_8 = pp_16_50;
  assign pp_0_51_0 = not_pp_9_51;
  assign pp_0_51_1 = pp_10_51;
  assign pp_0_51_2 = pp_11_51;
  assign pp_0_51_3 = pp_12_51;
  assign pp_0_51_4 = pp_13_51;
  assign pp_0_51_5 = pp_14_51;
  assign pp_0_51_6 = pp_15_51;
  assign pp_0_51_7 = pp_16_51;
  assign pp_0_52_0 = one;
  assign pp_0_52_1 = pp_10_52;
  assign pp_0_52_2 = pp_11_52;
  assign pp_0_52_3 = pp_12_52;
  assign pp_0_52_4 = pp_13_52;
  assign pp_0_52_5 = pp_14_52;
  assign pp_0_52_6 = pp_15_52;
  assign pp_0_52_7 = pp_16_52;
  assign pp_0_53_0 = not_pp_10_53;
  assign pp_0_53_1 = pp_11_53;
  assign pp_0_53_2 = pp_12_53;
  assign pp_0_53_3 = pp_13_53;
  assign pp_0_53_4 = pp_14_53;
  assign pp_0_53_5 = pp_15_53;
  assign pp_0_53_6 = pp_16_53;
  assign pp_0_54_0 = one;
  assign pp_0_54_1 = pp_11_54;
  assign pp_0_54_2 = pp_12_54;
  assign pp_0_54_3 = pp_13_54;
  assign pp_0_54_4 = pp_14_54;
  assign pp_0_54_5 = pp_15_54;
  assign pp_0_54_6 = pp_16_54;
  assign pp_0_55_0 = not_pp_11_55;
  assign pp_0_55_1 = pp_12_55;
  assign pp_0_55_2 = pp_13_55;
  assign pp_0_55_3 = pp_14_55;
  assign pp_0_55_4 = pp_15_55;
  assign pp_0_55_5 = pp_16_55;
  assign pp_0_56_0 = one;
  assign pp_0_56_1 = pp_12_56;
  assign pp_0_56_2 = pp_13_56;
  assign pp_0_56_3 = pp_14_56;
  assign pp_0_56_4 = pp_15_56;
  assign pp_0_56_5 = pp_16_56;
  assign pp_0_57_0 = not_pp_12_57;
  assign pp_0_57_1 = pp_13_57;
  assign pp_0_57_2 = pp_14_57;
  assign pp_0_57_3 = pp_15_57;
  assign pp_0_57_4 = pp_16_57;
  assign pp_0_58_0 = one;
  assign pp_0_58_1 = pp_13_58;
  assign pp_0_58_2 = pp_14_58;
  assign pp_0_58_3 = pp_15_58;
  assign pp_0_58_4 = pp_16_58;
  assign pp_0_59_0 = not_pp_13_59;
  assign pp_0_59_1 = pp_14_59;
  assign pp_0_59_2 = pp_15_59;
  assign pp_0_59_3 = pp_16_59;
  assign pp_0_60_0 = one;
  assign pp_0_60_1 = pp_14_60;
  assign pp_0_60_2 = pp_15_60;
  assign pp_0_60_3 = pp_16_60;
  assign pp_0_61_0 = not_pp_14_61;
  assign pp_0_61_1 = pp_15_61;
  assign pp_0_61_2 = pp_16_61;
  assign pp_0_62_0 = one;
  assign pp_0_62_1 = pp_15_62;
  assign pp_0_62_2 = pp_16_62;
  assign pp_0_63_0 = not_pp_15_63;
  assign pp_0_63_1 = pp_16_63;

  assign pp_1_0_0 = pp_0_0_0;
  assign pp_1_0_1 = pp_0_0_1;
  assign pp_1_1_0 = pp_0_1_0;
  MG_HA ha_0_2_0(
    .a(pp_0_2_0),
    .b(pp_0_2_1),
    .sum(pp_1_2_0),
    .cout(pp_1_3_0)
  );

  assign pp_1_2_1 = pp_0_2_2;
  MG_HA ha_0_3_0(
    .a(pp_0_3_0),
    .b(pp_0_3_1),
    .sum(pp_1_3_1),
    .cout(pp_1_4_0)
  );

  assign pp_1_4_1 = pp_0_4_0;
  assign pp_1_4_2 = pp_0_4_1;
  assign pp_1_4_3 = pp_0_4_2;
  assign pp_1_4_4 = pp_0_4_3;
  assign pp_1_5_0 = pp_0_5_0;
  assign pp_1_5_1 = pp_0_5_1;
  assign pp_1_5_2 = pp_0_5_2;
  MG_FA fa_0_6_0(
    .a(pp_0_6_0),
    .b(pp_0_6_1),
    .cin(pp_0_6_2),
    .sum(pp_1_6_0),
    .cout(pp_1_7_0)
  );

  assign pp_1_6_1 = pp_0_6_3;
  assign pp_1_6_2 = pp_0_6_4;
  MG_FA fa_0_7_0(
    .a(pp_0_7_0),
    .b(pp_0_7_1),
    .cin(pp_0_7_2),
    .sum(pp_1_7_1),
    .cout(pp_1_8_0)
  );

  assign pp_1_7_2 = pp_0_7_3;
  MG_FA fa_0_8_0(
    .a(pp_0_8_0),
    .b(pp_0_8_1),
    .cin(pp_0_8_2),
    .sum(pp_1_8_1),
    .cout(pp_1_9_0)
  );

  MG_FA fa_0_8_1(
    .a(pp_0_8_3),
    .b(pp_0_8_4),
    .cin(pp_0_8_5),
    .sum(pp_1_8_2),
    .cout(pp_1_9_1)
  );

  assign pp_1_9_2 = pp_0_9_0;
  assign pp_1_9_3 = pp_0_9_1;
  assign pp_1_9_4 = pp_0_9_2;
  assign pp_1_9_5 = pp_0_9_3;
  assign pp_1_9_6 = pp_0_9_4;
  MG_FA fa_0_10_0(
    .a(pp_0_10_0),
    .b(pp_0_10_1),
    .cin(pp_0_10_2),
    .sum(pp_1_10_0),
    .cout(pp_1_11_0)
  );

  MG_FA fa_0_10_1(
    .a(pp_0_10_3),
    .b(pp_0_10_4),
    .cin(pp_0_10_5),
    .sum(pp_1_10_1),
    .cout(pp_1_11_1)
  );

  assign pp_1_10_2 = pp_0_10_6;
  MG_FA fa_0_11_0(
    .a(pp_0_11_0),
    .b(pp_0_11_1),
    .cin(pp_0_11_2),
    .sum(pp_1_11_2),
    .cout(pp_1_12_0)
  );

  MG_FA fa_0_11_1(
    .a(pp_0_11_3),
    .b(pp_0_11_4),
    .cin(pp_0_11_5),
    .sum(pp_1_11_3),
    .cout(pp_1_12_1)
  );

  MG_FA fa_0_12_0(
    .a(pp_0_12_0),
    .b(pp_0_12_1),
    .cin(pp_0_12_2),
    .sum(pp_1_12_2),
    .cout(pp_1_13_0)
  );

  MG_FA fa_0_12_1(
    .a(pp_0_12_3),
    .b(pp_0_12_4),
    .cin(pp_0_12_5),
    .sum(pp_1_12_3),
    .cout(pp_1_13_1)
  );

  assign pp_1_12_4 = pp_0_12_6;
  assign pp_1_12_5 = pp_0_12_7;
  MG_FA fa_0_13_0(
    .a(pp_0_13_0),
    .b(pp_0_13_1),
    .cin(pp_0_13_2),
    .sum(pp_1_13_2),
    .cout(pp_1_14_0)
  );

  assign pp_1_13_3 = pp_0_13_3;
  assign pp_1_13_4 = pp_0_13_4;
  assign pp_1_13_5 = pp_0_13_5;
  assign pp_1_13_6 = pp_0_13_6;
  MG_FA fa_0_14_0(
    .a(pp_0_14_0),
    .b(pp_0_14_1),
    .cin(pp_0_14_2),
    .sum(pp_1_14_1),
    .cout(pp_1_15_0)
  );

  MG_FA fa_0_14_1(
    .a(pp_0_14_3),
    .b(pp_0_14_4),
    .cin(pp_0_14_5),
    .sum(pp_1_14_2),
    .cout(pp_1_15_1)
  );

  MG_FA fa_0_14_2(
    .a(pp_0_14_6),
    .b(pp_0_14_7),
    .cin(pp_0_14_8),
    .sum(pp_1_14_3),
    .cout(pp_1_15_2)
  );

  MG_FA fa_0_15_0(
    .a(pp_0_15_0),
    .b(pp_0_15_1),
    .cin(pp_0_15_2),
    .sum(pp_1_15_3),
    .cout(pp_1_16_0)
  );

  MG_FA fa_0_15_1(
    .a(pp_0_15_3),
    .b(pp_0_15_4),
    .cin(pp_0_15_5),
    .sum(pp_1_15_4),
    .cout(pp_1_16_1)
  );

  assign pp_1_15_5 = pp_0_15_6;
  assign pp_1_15_6 = pp_0_15_7;
  MG_FA fa_0_16_0(
    .a(pp_0_16_0),
    .b(pp_0_16_1),
    .cin(pp_0_16_2),
    .sum(pp_1_16_2),
    .cout(pp_1_17_0)
  );

  MG_FA fa_0_16_1(
    .a(pp_0_16_3),
    .b(pp_0_16_4),
    .cin(pp_0_16_5),
    .sum(pp_1_16_3),
    .cout(pp_1_17_1)
  );

  MG_FA fa_0_16_2(
    .a(pp_0_16_6),
    .b(pp_0_16_7),
    .cin(pp_0_16_8),
    .sum(pp_1_16_4),
    .cout(pp_1_17_2)
  );

  assign pp_1_16_5 = pp_0_16_9;
  MG_FA fa_0_17_0(
    .a(pp_0_17_0),
    .b(pp_0_17_1),
    .cin(pp_0_17_2),
    .sum(pp_1_17_3),
    .cout(pp_1_18_0)
  );

  MG_FA fa_0_17_1(
    .a(pp_0_17_3),
    .b(pp_0_17_4),
    .cin(pp_0_17_5),
    .sum(pp_1_17_4),
    .cout(pp_1_18_1)
  );

  MG_FA fa_0_17_2(
    .a(pp_0_17_6),
    .b(pp_0_17_7),
    .cin(pp_0_17_8),
    .sum(pp_1_17_5),
    .cout(pp_1_18_2)
  );

  MG_FA fa_0_18_0(
    .a(pp_0_18_0),
    .b(pp_0_18_1),
    .cin(pp_0_18_2),
    .sum(pp_1_18_3),
    .cout(pp_1_19_0)
  );

  MG_FA fa_0_18_1(
    .a(pp_0_18_3),
    .b(pp_0_18_4),
    .cin(pp_0_18_5),
    .sum(pp_1_18_4),
    .cout(pp_1_19_1)
  );

  assign pp_1_18_5 = pp_0_18_6;
  assign pp_1_18_6 = pp_0_18_7;
  assign pp_1_18_7 = pp_0_18_8;
  assign pp_1_18_8 = pp_0_18_9;
  assign pp_1_18_9 = pp_0_18_10;
  MG_FA fa_0_19_0(
    .a(pp_0_19_0),
    .b(pp_0_19_1),
    .cin(pp_0_19_2),
    .sum(pp_1_19_2),
    .cout(pp_1_20_0)
  );

  MG_FA fa_0_19_1(
    .a(pp_0_19_3),
    .b(pp_0_19_4),
    .cin(pp_0_19_5),
    .sum(pp_1_19_3),
    .cout(pp_1_20_1)
  );

  MG_FA fa_0_19_2(
    .a(pp_0_19_6),
    .b(pp_0_19_7),
    .cin(pp_0_19_8),
    .sum(pp_1_19_4),
    .cout(pp_1_20_2)
  );

  assign pp_1_19_5 = pp_0_19_9;
  MG_FA fa_0_20_0(
    .a(pp_0_20_0),
    .b(pp_0_20_1),
    .cin(pp_0_20_2),
    .sum(pp_1_20_3),
    .cout(pp_1_21_0)
  );

  MG_FA fa_0_20_1(
    .a(pp_0_20_3),
    .b(pp_0_20_4),
    .cin(pp_0_20_5),
    .sum(pp_1_20_4),
    .cout(pp_1_21_1)
  );

  MG_FA fa_0_20_2(
    .a(pp_0_20_6),
    .b(pp_0_20_7),
    .cin(pp_0_20_8),
    .sum(pp_1_20_5),
    .cout(pp_1_21_2)
  );

  MG_FA fa_0_20_3(
    .a(pp_0_20_9),
    .b(pp_0_20_10),
    .cin(pp_0_20_11),
    .sum(pp_1_20_6),
    .cout(pp_1_21_3)
  );

  MG_FA fa_0_21_0(
    .a(pp_0_21_0),
    .b(pp_0_21_1),
    .cin(pp_0_21_2),
    .sum(pp_1_21_4),
    .cout(pp_1_22_0)
  );

  MG_FA fa_0_21_1(
    .a(pp_0_21_3),
    .b(pp_0_21_4),
    .cin(pp_0_21_5),
    .sum(pp_1_21_5),
    .cout(pp_1_22_1)
  );

  MG_FA fa_0_21_2(
    .a(pp_0_21_6),
    .b(pp_0_21_7),
    .cin(pp_0_21_8),
    .sum(pp_1_21_6),
    .cout(pp_1_22_2)
  );

  assign pp_1_21_7 = pp_0_21_9;
  assign pp_1_21_8 = pp_0_21_10;
  MG_FA fa_0_22_0(
    .a(pp_0_22_0),
    .b(pp_0_22_1),
    .cin(pp_0_22_2),
    .sum(pp_1_22_3),
    .cout(pp_1_23_0)
  );

  MG_FA fa_0_22_1(
    .a(pp_0_22_3),
    .b(pp_0_22_4),
    .cin(pp_0_22_5),
    .sum(pp_1_22_4),
    .cout(pp_1_23_1)
  );

  MG_FA fa_0_22_2(
    .a(pp_0_22_6),
    .b(pp_0_22_7),
    .cin(pp_0_22_8),
    .sum(pp_1_22_5),
    .cout(pp_1_23_2)
  );

  MG_FA fa_0_22_3(
    .a(pp_0_22_9),
    .b(pp_0_22_10),
    .cin(pp_0_22_11),
    .sum(pp_1_22_6),
    .cout(pp_1_23_3)
  );

  assign pp_1_22_7 = pp_0_22_12;
  MG_FA fa_0_23_0(
    .a(pp_0_23_0),
    .b(pp_0_23_1),
    .cin(pp_0_23_2),
    .sum(pp_1_23_4),
    .cout(pp_1_24_0)
  );

  MG_FA fa_0_23_1(
    .a(pp_0_23_3),
    .b(pp_0_23_4),
    .cin(pp_0_23_5),
    .sum(pp_1_23_5),
    .cout(pp_1_24_1)
  );

  MG_FA fa_0_23_2(
    .a(pp_0_23_6),
    .b(pp_0_23_7),
    .cin(pp_0_23_8),
    .sum(pp_1_23_6),
    .cout(pp_1_24_2)
  );

  MG_FA fa_0_23_3(
    .a(pp_0_23_9),
    .b(pp_0_23_10),
    .cin(pp_0_23_11),
    .sum(pp_1_23_7),
    .cout(pp_1_24_3)
  );

  MG_FA fa_0_24_0(
    .a(pp_0_24_0),
    .b(pp_0_24_1),
    .cin(pp_0_24_2),
    .sum(pp_1_24_4),
    .cout(pp_1_25_0)
  );

  MG_FA fa_0_24_1(
    .a(pp_0_24_3),
    .b(pp_0_24_4),
    .cin(pp_0_24_5),
    .sum(pp_1_24_5),
    .cout(pp_1_25_1)
  );

  MG_FA fa_0_24_2(
    .a(pp_0_24_6),
    .b(pp_0_24_7),
    .cin(pp_0_24_8),
    .sum(pp_1_24_6),
    .cout(pp_1_25_2)
  );

  MG_FA fa_0_24_3(
    .a(pp_0_24_9),
    .b(pp_0_24_10),
    .cin(pp_0_24_11),
    .sum(pp_1_24_7),
    .cout(pp_1_25_3)
  );

  assign pp_1_24_8 = pp_0_24_12;
  assign pp_1_24_9 = pp_0_24_13;
  MG_FA fa_0_25_0(
    .a(pp_0_25_0),
    .b(pp_0_25_1),
    .cin(pp_0_25_2),
    .sum(pp_1_25_4),
    .cout(pp_1_26_0)
  );

  MG_FA fa_0_25_1(
    .a(pp_0_25_3),
    .b(pp_0_25_4),
    .cin(pp_0_25_5),
    .sum(pp_1_25_5),
    .cout(pp_1_26_1)
  );

  MG_FA fa_0_25_2(
    .a(pp_0_25_6),
    .b(pp_0_25_7),
    .cin(pp_0_25_8),
    .sum(pp_1_25_6),
    .cout(pp_1_26_2)
  );

  MG_FA fa_0_25_3(
    .a(pp_0_25_9),
    .b(pp_0_25_10),
    .cin(pp_0_25_11),
    .sum(pp_1_25_7),
    .cout(pp_1_26_3)
  );

  assign pp_1_25_8 = pp_0_25_12;
  MG_FA fa_0_26_0(
    .a(pp_0_26_0),
    .b(pp_0_26_1),
    .cin(pp_0_26_2),
    .sum(pp_1_26_4),
    .cout(pp_1_27_0)
  );

  MG_FA fa_0_26_1(
    .a(pp_0_26_3),
    .b(pp_0_26_4),
    .cin(pp_0_26_5),
    .sum(pp_1_26_5),
    .cout(pp_1_27_1)
  );

  MG_FA fa_0_26_2(
    .a(pp_0_26_6),
    .b(pp_0_26_7),
    .cin(pp_0_26_8),
    .sum(pp_1_26_6),
    .cout(pp_1_27_2)
  );

  MG_FA fa_0_26_3(
    .a(pp_0_26_9),
    .b(pp_0_26_10),
    .cin(pp_0_26_11),
    .sum(pp_1_26_7),
    .cout(pp_1_27_3)
  );

  MG_FA fa_0_26_4(
    .a(pp_0_26_12),
    .b(pp_0_26_13),
    .cin(pp_0_26_14),
    .sum(pp_1_26_8),
    .cout(pp_1_27_4)
  );

  MG_FA fa_0_27_0(
    .a(pp_0_27_0),
    .b(pp_0_27_1),
    .cin(pp_0_27_2),
    .sum(pp_1_27_5),
    .cout(pp_1_28_0)
  );

  MG_FA fa_0_27_1(
    .a(pp_0_27_3),
    .b(pp_0_27_4),
    .cin(pp_0_27_5),
    .sum(pp_1_27_6),
    .cout(pp_1_28_1)
  );

  MG_FA fa_0_27_2(
    .a(pp_0_27_6),
    .b(pp_0_27_7),
    .cin(pp_0_27_8),
    .sum(pp_1_27_7),
    .cout(pp_1_28_2)
  );

  assign pp_1_27_8 = pp_0_27_9;
  assign pp_1_27_9 = pp_0_27_10;
  assign pp_1_27_10 = pp_0_27_11;
  assign pp_1_27_11 = pp_0_27_12;
  assign pp_1_27_12 = pp_0_27_13;
  MG_FA fa_0_28_0(
    .a(pp_0_28_0),
    .b(pp_0_28_1),
    .cin(pp_0_28_2),
    .sum(pp_1_28_3),
    .cout(pp_1_29_0)
  );

  MG_FA fa_0_28_1(
    .a(pp_0_28_3),
    .b(pp_0_28_4),
    .cin(pp_0_28_5),
    .sum(pp_1_28_4),
    .cout(pp_1_29_1)
  );

  MG_FA fa_0_28_2(
    .a(pp_0_28_6),
    .b(pp_0_28_7),
    .cin(pp_0_28_8),
    .sum(pp_1_28_5),
    .cout(pp_1_29_2)
  );

  MG_FA fa_0_28_3(
    .a(pp_0_28_9),
    .b(pp_0_28_10),
    .cin(pp_0_28_11),
    .sum(pp_1_28_6),
    .cout(pp_1_29_3)
  );

  MG_FA fa_0_28_4(
    .a(pp_0_28_12),
    .b(pp_0_28_13),
    .cin(pp_0_28_14),
    .sum(pp_1_28_7),
    .cout(pp_1_29_4)
  );

  assign pp_1_28_8 = pp_0_28_15;
  MG_FA fa_0_29_0(
    .a(pp_0_29_0),
    .b(pp_0_29_1),
    .cin(pp_0_29_2),
    .sum(pp_1_29_5),
    .cout(pp_1_30_0)
  );

  MG_FA fa_0_29_1(
    .a(pp_0_29_3),
    .b(pp_0_29_4),
    .cin(pp_0_29_5),
    .sum(pp_1_29_6),
    .cout(pp_1_30_1)
  );

  MG_FA fa_0_29_2(
    .a(pp_0_29_6),
    .b(pp_0_29_7),
    .cin(pp_0_29_8),
    .sum(pp_1_29_7),
    .cout(pp_1_30_2)
  );

  MG_FA fa_0_29_3(
    .a(pp_0_29_9),
    .b(pp_0_29_10),
    .cin(pp_0_29_11),
    .sum(pp_1_29_8),
    .cout(pp_1_30_3)
  );

  MG_FA fa_0_29_4(
    .a(pp_0_29_12),
    .b(pp_0_29_13),
    .cin(pp_0_29_14),
    .sum(pp_1_29_9),
    .cout(pp_1_30_4)
  );

  MG_FA fa_0_30_0(
    .a(pp_0_30_0),
    .b(pp_0_30_1),
    .cin(pp_0_30_2),
    .sum(pp_1_30_5),
    .cout(pp_1_31_0)
  );

  MG_FA fa_0_30_1(
    .a(pp_0_30_3),
    .b(pp_0_30_4),
    .cin(pp_0_30_5),
    .sum(pp_1_30_6),
    .cout(pp_1_31_1)
  );

  MG_FA fa_0_30_2(
    .a(pp_0_30_6),
    .b(pp_0_30_7),
    .cin(pp_0_30_8),
    .sum(pp_1_30_7),
    .cout(pp_1_31_2)
  );

  MG_FA fa_0_30_3(
    .a(pp_0_30_9),
    .b(pp_0_30_10),
    .cin(pp_0_30_11),
    .sum(pp_1_30_8),
    .cout(pp_1_31_3)
  );

  MG_FA fa_0_30_4(
    .a(pp_0_30_12),
    .b(pp_0_30_13),
    .cin(pp_0_30_14),
    .sum(pp_1_30_9),
    .cout(pp_1_31_4)
  );

  assign pp_1_30_10 = pp_0_30_15;
  assign pp_1_30_11 = pp_0_30_16;
  MG_FA fa_0_31_0(
    .a(pp_0_31_0),
    .b(pp_0_31_1),
    .cin(pp_0_31_2),
    .sum(pp_1_31_5),
    .cout(pp_1_32_0)
  );

  MG_FA fa_0_31_1(
    .a(pp_0_31_3),
    .b(pp_0_31_4),
    .cin(pp_0_31_5),
    .sum(pp_1_31_6),
    .cout(pp_1_32_1)
  );

  MG_FA fa_0_31_2(
    .a(pp_0_31_6),
    .b(pp_0_31_7),
    .cin(pp_0_31_8),
    .sum(pp_1_31_7),
    .cout(pp_1_32_2)
  );

  MG_FA fa_0_31_3(
    .a(pp_0_31_9),
    .b(pp_0_31_10),
    .cin(pp_0_31_11),
    .sum(pp_1_31_8),
    .cout(pp_1_32_3)
  );

  MG_HA ha_0_31_4(
    .a(pp_0_31_12),
    .b(pp_0_31_13),
    .sum(pp_1_31_9),
    .cout(pp_1_32_4)
  );

  assign pp_1_31_10 = pp_0_31_14;
  assign pp_1_31_11 = pp_0_31_15;
  MG_FA fa_0_32_0(
    .a(pp_0_32_0),
    .b(pp_0_32_1),
    .cin(pp_0_32_2),
    .sum(pp_1_32_5),
    .cout(pp_1_33_0)
  );

  MG_FA fa_0_32_1(
    .a(pp_0_32_3),
    .b(pp_0_32_4),
    .cin(pp_0_32_5),
    .sum(pp_1_32_6),
    .cout(pp_1_33_1)
  );

  MG_FA fa_0_32_2(
    .a(pp_0_32_6),
    .b(pp_0_32_7),
    .cin(pp_0_32_8),
    .sum(pp_1_32_7),
    .cout(pp_1_33_2)
  );

  MG_FA fa_0_32_3(
    .a(pp_0_32_9),
    .b(pp_0_32_10),
    .cin(pp_0_32_11),
    .sum(pp_1_32_8),
    .cout(pp_1_33_3)
  );

  MG_FA fa_0_32_4(
    .a(pp_0_32_12),
    .b(pp_0_32_13),
    .cin(pp_0_32_14),
    .sum(pp_1_32_9),
    .cout(pp_1_33_4)
  );

  assign pp_1_32_10 = pp_0_32_15;
  assign pp_1_32_11 = pp_0_32_16;
  MG_FA fa_0_33_0(
    .a(pp_0_33_0),
    .b(pp_0_33_1),
    .cin(pp_0_33_2),
    .sum(pp_1_33_5),
    .cout(pp_1_34_0)
  );

  MG_FA fa_0_33_1(
    .a(pp_0_33_3),
    .b(pp_0_33_4),
    .cin(pp_0_33_5),
    .sum(pp_1_33_6),
    .cout(pp_1_34_1)
  );

  MG_FA fa_0_33_2(
    .a(pp_0_33_6),
    .b(pp_0_33_7),
    .cin(pp_0_33_8),
    .sum(pp_1_33_7),
    .cout(pp_1_34_2)
  );

  MG_FA fa_0_33_3(
    .a(pp_0_33_9),
    .b(pp_0_33_10),
    .cin(pp_0_33_11),
    .sum(pp_1_33_8),
    .cout(pp_1_34_3)
  );

  MG_FA fa_0_33_4(
    .a(pp_0_33_12),
    .b(pp_0_33_13),
    .cin(pp_0_33_14),
    .sum(pp_1_33_9),
    .cout(pp_1_34_4)
  );

  assign pp_1_33_10 = pp_0_33_15;
  assign pp_1_33_11 = pp_0_33_16;
  MG_FA fa_0_34_0(
    .a(pp_0_34_0),
    .b(pp_0_34_1),
    .cin(pp_0_34_2),
    .sum(pp_1_34_5),
    .cout(pp_1_35_0)
  );

  MG_FA fa_0_34_1(
    .a(pp_0_34_3),
    .b(pp_0_34_4),
    .cin(pp_0_34_5),
    .sum(pp_1_34_6),
    .cout(pp_1_35_1)
  );

  MG_FA fa_0_34_2(
    .a(pp_0_34_6),
    .b(pp_0_34_7),
    .cin(pp_0_34_8),
    .sum(pp_1_34_7),
    .cout(pp_1_35_2)
  );

  MG_FA fa_0_34_3(
    .a(pp_0_34_9),
    .b(pp_0_34_10),
    .cin(pp_0_34_11),
    .sum(pp_1_34_8),
    .cout(pp_1_35_3)
  );

  MG_FA fa_0_34_4(
    .a(pp_0_34_12),
    .b(pp_0_34_13),
    .cin(pp_0_34_14),
    .sum(pp_1_34_9),
    .cout(pp_1_35_4)
  );

  assign pp_1_34_10 = pp_0_34_15;
  assign pp_1_34_11 = pp_0_34_16;
  MG_FA fa_0_35_0(
    .a(pp_0_35_0),
    .b(pp_0_35_1),
    .cin(pp_0_35_2),
    .sum(pp_1_35_5),
    .cout(pp_1_36_0)
  );

  MG_FA fa_0_35_1(
    .a(pp_0_35_3),
    .b(pp_0_35_4),
    .cin(pp_0_35_5),
    .sum(pp_1_35_6),
    .cout(pp_1_36_1)
  );

  MG_FA fa_0_35_2(
    .a(pp_0_35_6),
    .b(pp_0_35_7),
    .cin(pp_0_35_8),
    .sum(pp_1_35_7),
    .cout(pp_1_36_2)
  );

  MG_FA fa_0_35_3(
    .a(pp_0_35_9),
    .b(pp_0_35_10),
    .cin(pp_0_35_11),
    .sum(pp_1_35_8),
    .cout(pp_1_36_3)
  );

  MG_FA fa_0_35_4(
    .a(pp_0_35_12),
    .b(pp_0_35_13),
    .cin(pp_0_35_14),
    .sum(pp_1_35_9),
    .cout(pp_1_36_4)
  );

  assign pp_1_35_10 = pp_0_35_15;
  assign pp_1_35_11 = pp_0_35_16;
  MG_FA fa_0_36_0(
    .a(pp_0_36_0),
    .b(pp_0_36_1),
    .cin(pp_0_36_2),
    .sum(pp_1_36_5),
    .cout(pp_1_37_0)
  );

  MG_FA fa_0_36_1(
    .a(pp_0_36_3),
    .b(pp_0_36_4),
    .cin(pp_0_36_5),
    .sum(pp_1_36_6),
    .cout(pp_1_37_1)
  );

  MG_FA fa_0_36_2(
    .a(pp_0_36_6),
    .b(pp_0_36_7),
    .cin(pp_0_36_8),
    .sum(pp_1_36_7),
    .cout(pp_1_37_2)
  );

  MG_FA fa_0_36_3(
    .a(pp_0_36_9),
    .b(pp_0_36_10),
    .cin(pp_0_36_11),
    .sum(pp_1_36_8),
    .cout(pp_1_37_3)
  );

  MG_FA fa_0_36_4(
    .a(pp_0_36_12),
    .b(pp_0_36_13),
    .cin(pp_0_36_14),
    .sum(pp_1_36_9),
    .cout(pp_1_37_4)
  );

  assign pp_1_36_10 = pp_0_36_15;
  MG_FA fa_0_37_0(
    .a(pp_0_37_0),
    .b(pp_0_37_1),
    .cin(pp_0_37_2),
    .sum(pp_1_37_5),
    .cout(pp_1_38_0)
  );

  MG_FA fa_0_37_1(
    .a(pp_0_37_3),
    .b(pp_0_37_4),
    .cin(pp_0_37_5),
    .sum(pp_1_37_6),
    .cout(pp_1_38_1)
  );

  MG_FA fa_0_37_2(
    .a(pp_0_37_6),
    .b(pp_0_37_7),
    .cin(pp_0_37_8),
    .sum(pp_1_37_7),
    .cout(pp_1_38_2)
  );

  MG_FA fa_0_37_3(
    .a(pp_0_37_9),
    .b(pp_0_37_10),
    .cin(pp_0_37_11),
    .sum(pp_1_37_8),
    .cout(pp_1_38_3)
  );

  assign pp_1_37_9 = pp_0_37_12;
  assign pp_1_37_10 = pp_0_37_13;
  assign pp_1_37_11 = pp_0_37_14;
  MG_FA fa_0_38_0(
    .a(pp_0_38_0),
    .b(pp_0_38_1),
    .cin(pp_0_38_2),
    .sum(pp_1_38_4),
    .cout(pp_1_39_0)
  );

  MG_FA fa_0_38_1(
    .a(pp_0_38_3),
    .b(pp_0_38_4),
    .cin(pp_0_38_5),
    .sum(pp_1_38_5),
    .cout(pp_1_39_1)
  );

  MG_FA fa_0_38_2(
    .a(pp_0_38_6),
    .b(pp_0_38_7),
    .cin(pp_0_38_8),
    .sum(pp_1_38_6),
    .cout(pp_1_39_2)
  );

  MG_FA fa_0_38_3(
    .a(pp_0_38_9),
    .b(pp_0_38_10),
    .cin(pp_0_38_11),
    .sum(pp_1_38_7),
    .cout(pp_1_39_3)
  );

  MG_FA fa_0_38_4(
    .a(pp_0_38_12),
    .b(pp_0_38_13),
    .cin(pp_0_38_14),
    .sum(pp_1_38_8),
    .cout(pp_1_39_4)
  );

  MG_FA fa_0_39_0(
    .a(pp_0_39_0),
    .b(pp_0_39_1),
    .cin(pp_0_39_2),
    .sum(pp_1_39_5),
    .cout(pp_1_40_0)
  );

  MG_FA fa_0_39_1(
    .a(pp_0_39_3),
    .b(pp_0_39_4),
    .cin(pp_0_39_5),
    .sum(pp_1_39_6),
    .cout(pp_1_40_1)
  );

  MG_FA fa_0_39_2(
    .a(pp_0_39_6),
    .b(pp_0_39_7),
    .cin(pp_0_39_8),
    .sum(pp_1_39_7),
    .cout(pp_1_40_2)
  );

  MG_FA fa_0_39_3(
    .a(pp_0_39_9),
    .b(pp_0_39_10),
    .cin(pp_0_39_11),
    .sum(pp_1_39_8),
    .cout(pp_1_40_3)
  );

  assign pp_1_39_9 = pp_0_39_12;
  assign pp_1_39_10 = pp_0_39_13;
  MG_FA fa_0_40_0(
    .a(pp_0_40_0),
    .b(pp_0_40_1),
    .cin(pp_0_40_2),
    .sum(pp_1_40_4),
    .cout(pp_1_41_0)
  );

  MG_FA fa_0_40_1(
    .a(pp_0_40_3),
    .b(pp_0_40_4),
    .cin(pp_0_40_5),
    .sum(pp_1_40_5),
    .cout(pp_1_41_1)
  );

  MG_FA fa_0_40_2(
    .a(pp_0_40_6),
    .b(pp_0_40_7),
    .cin(pp_0_40_8),
    .sum(pp_1_40_6),
    .cout(pp_1_41_2)
  );

  MG_FA fa_0_40_3(
    .a(pp_0_40_9),
    .b(pp_0_40_10),
    .cin(pp_0_40_11),
    .sum(pp_1_40_7),
    .cout(pp_1_41_3)
  );

  assign pp_1_40_8 = pp_0_40_12;
  assign pp_1_40_9 = pp_0_40_13;
  MG_FA fa_0_41_0(
    .a(pp_0_41_0),
    .b(pp_0_41_1),
    .cin(pp_0_41_2),
    .sum(pp_1_41_4),
    .cout(pp_1_42_0)
  );

  MG_FA fa_0_41_1(
    .a(pp_0_41_3),
    .b(pp_0_41_4),
    .cin(pp_0_41_5),
    .sum(pp_1_41_5),
    .cout(pp_1_42_1)
  );

  MG_FA fa_0_41_2(
    .a(pp_0_41_6),
    .b(pp_0_41_7),
    .cin(pp_0_41_8),
    .sum(pp_1_41_6),
    .cout(pp_1_42_2)
  );

  MG_FA fa_0_41_3(
    .a(pp_0_41_9),
    .b(pp_0_41_10),
    .cin(pp_0_41_11),
    .sum(pp_1_41_7),
    .cout(pp_1_42_3)
  );

  assign pp_1_41_8 = pp_0_41_12;
  MG_FA fa_0_42_0(
    .a(pp_0_42_0),
    .b(pp_0_42_1),
    .cin(pp_0_42_2),
    .sum(pp_1_42_4),
    .cout(pp_1_43_0)
  );

  MG_FA fa_0_42_1(
    .a(pp_0_42_3),
    .b(pp_0_42_4),
    .cin(pp_0_42_5),
    .sum(pp_1_42_5),
    .cout(pp_1_43_1)
  );

  MG_FA fa_0_42_2(
    .a(pp_0_42_6),
    .b(pp_0_42_7),
    .cin(pp_0_42_8),
    .sum(pp_1_42_6),
    .cout(pp_1_43_2)
  );

  MG_FA fa_0_42_3(
    .a(pp_0_42_9),
    .b(pp_0_42_10),
    .cin(pp_0_42_11),
    .sum(pp_1_42_7),
    .cout(pp_1_43_3)
  );

  assign pp_1_42_8 = pp_0_42_12;
  MG_FA fa_0_43_0(
    .a(pp_0_43_0),
    .b(pp_0_43_1),
    .cin(pp_0_43_2),
    .sum(pp_1_43_4),
    .cout(pp_1_44_0)
  );

  MG_FA fa_0_43_1(
    .a(pp_0_43_3),
    .b(pp_0_43_4),
    .cin(pp_0_43_5),
    .sum(pp_1_43_5),
    .cout(pp_1_44_1)
  );

  assign pp_1_43_6 = pp_0_43_6;
  assign pp_1_43_7 = pp_0_43_7;
  assign pp_1_43_8 = pp_0_43_8;
  assign pp_1_43_9 = pp_0_43_9;
  assign pp_1_43_10 = pp_0_43_10;
  assign pp_1_43_11 = pp_0_43_11;
  MG_FA fa_0_44_0(
    .a(pp_0_44_0),
    .b(pp_0_44_1),
    .cin(pp_0_44_2),
    .sum(pp_1_44_2),
    .cout(pp_1_45_0)
  );

  MG_FA fa_0_44_1(
    .a(pp_0_44_3),
    .b(pp_0_44_4),
    .cin(pp_0_44_5),
    .sum(pp_1_44_3),
    .cout(pp_1_45_1)
  );

  MG_FA fa_0_44_2(
    .a(pp_0_44_6),
    .b(pp_0_44_7),
    .cin(pp_0_44_8),
    .sum(pp_1_44_4),
    .cout(pp_1_45_2)
  );

  MG_FA fa_0_44_3(
    .a(pp_0_44_9),
    .b(pp_0_44_10),
    .cin(pp_0_44_11),
    .sum(pp_1_44_5),
    .cout(pp_1_45_3)
  );

  MG_FA fa_0_45_0(
    .a(pp_0_45_0),
    .b(pp_0_45_1),
    .cin(pp_0_45_2),
    .sum(pp_1_45_4),
    .cout(pp_1_46_0)
  );

  assign pp_1_45_5 = pp_0_45_3;
  assign pp_1_45_6 = pp_0_45_4;
  assign pp_1_45_7 = pp_0_45_5;
  assign pp_1_45_8 = pp_0_45_6;
  assign pp_1_45_9 = pp_0_45_7;
  assign pp_1_45_10 = pp_0_45_8;
  assign pp_1_45_11 = pp_0_45_9;
  assign pp_1_45_12 = pp_0_45_10;
  MG_FA fa_0_46_0(
    .a(pp_0_46_0),
    .b(pp_0_46_1),
    .cin(pp_0_46_2),
    .sum(pp_1_46_1),
    .cout(pp_1_47_0)
  );

  MG_HA ha_0_46_1(
    .a(pp_0_46_3),
    .b(pp_0_46_4),
    .sum(pp_1_46_2),
    .cout(pp_1_47_1)
  );

  assign pp_1_46_3 = pp_0_46_5;
  assign pp_1_46_4 = pp_0_46_6;
  assign pp_1_46_5 = pp_0_46_7;
  assign pp_1_46_6 = pp_0_46_8;
  assign pp_1_46_7 = pp_0_46_9;
  assign pp_1_46_8 = pp_0_46_10;
  MG_FA fa_0_47_0(
    .a(pp_0_47_0),
    .b(pp_0_47_1),
    .cin(pp_0_47_2),
    .sum(pp_1_47_2),
    .cout(pp_1_48_0)
  );

  MG_FA fa_0_47_1(
    .a(pp_0_47_3),
    .b(pp_0_47_4),
    .cin(pp_0_47_5),
    .sum(pp_1_47_3),
    .cout(pp_1_48_1)
  );

  MG_FA fa_0_47_2(
    .a(pp_0_47_6),
    .b(pp_0_47_7),
    .cin(pp_0_47_8),
    .sum(pp_1_47_4),
    .cout(pp_1_48_2)
  );

  assign pp_1_47_5 = pp_0_47_9;
  MG_FA fa_0_48_0(
    .a(pp_0_48_0),
    .b(pp_0_48_1),
    .cin(pp_0_48_2),
    .sum(pp_1_48_3),
    .cout(pp_1_49_0)
  );

  MG_FA fa_0_48_1(
    .a(pp_0_48_3),
    .b(pp_0_48_4),
    .cin(pp_0_48_5),
    .sum(pp_1_48_4),
    .cout(pp_1_49_1)
  );

  assign pp_1_48_5 = pp_0_48_6;
  assign pp_1_48_6 = pp_0_48_7;
  assign pp_1_48_7 = pp_0_48_8;
  assign pp_1_48_8 = pp_0_48_9;
  MG_FA fa_0_49_0(
    .a(pp_0_49_0),
    .b(pp_0_49_1),
    .cin(pp_0_49_2),
    .sum(pp_1_49_2),
    .cout(pp_1_50_0)
  );

  MG_FA fa_0_49_1(
    .a(pp_0_49_3),
    .b(pp_0_49_4),
    .cin(pp_0_49_5),
    .sum(pp_1_49_3),
    .cout(pp_1_50_1)
  );

  MG_FA fa_0_49_2(
    .a(pp_0_49_6),
    .b(pp_0_49_7),
    .cin(pp_0_49_8),
    .sum(pp_1_49_4),
    .cout(pp_1_50_2)
  );

  MG_FA fa_0_50_0(
    .a(pp_0_50_0),
    .b(pp_0_50_1),
    .cin(pp_0_50_2),
    .sum(pp_1_50_3),
    .cout(pp_1_51_0)
  );

  MG_FA fa_0_50_1(
    .a(pp_0_50_3),
    .b(pp_0_50_4),
    .cin(pp_0_50_5),
    .sum(pp_1_50_4),
    .cout(pp_1_51_1)
  );

  MG_FA fa_0_50_2(
    .a(pp_0_50_6),
    .b(pp_0_50_7),
    .cin(pp_0_50_8),
    .sum(pp_1_50_5),
    .cout(pp_1_51_2)
  );

  MG_FA fa_0_51_0(
    .a(pp_0_51_0),
    .b(pp_0_51_1),
    .cin(pp_0_51_2),
    .sum(pp_1_51_3),
    .cout(pp_1_52_0)
  );

  MG_FA fa_0_51_1(
    .a(pp_0_51_3),
    .b(pp_0_51_4),
    .cin(pp_0_51_5),
    .sum(pp_1_51_4),
    .cout(pp_1_52_1)
  );

  assign pp_1_51_5 = pp_0_51_6;
  assign pp_1_51_6 = pp_0_51_7;
  MG_FA fa_0_52_0(
    .a(pp_0_52_0),
    .b(pp_0_52_1),
    .cin(pp_0_52_2),
    .sum(pp_1_52_2),
    .cout(pp_1_53_0)
  );

  MG_FA fa_0_52_1(
    .a(pp_0_52_3),
    .b(pp_0_52_4),
    .cin(pp_0_52_5),
    .sum(pp_1_52_3),
    .cout(pp_1_53_1)
  );

  assign pp_1_52_4 = pp_0_52_6;
  assign pp_1_52_5 = pp_0_52_7;
  assign pp_1_53_2 = pp_0_53_0;
  assign pp_1_53_3 = pp_0_53_1;
  assign pp_1_53_4 = pp_0_53_2;
  assign pp_1_53_5 = pp_0_53_3;
  assign pp_1_53_6 = pp_0_53_4;
  assign pp_1_53_7 = pp_0_53_5;
  assign pp_1_53_8 = pp_0_53_6;
  MG_FA fa_0_54_0(
    .a(pp_0_54_0),
    .b(pp_0_54_1),
    .cin(pp_0_54_2),
    .sum(pp_1_54_0),
    .cout(pp_1_55_0)
  );

  MG_FA fa_0_54_1(
    .a(pp_0_54_3),
    .b(pp_0_54_4),
    .cin(pp_0_54_5),
    .sum(pp_1_54_1),
    .cout(pp_1_55_1)
  );

  assign pp_1_54_2 = pp_0_54_6;
  MG_FA fa_0_55_0(
    .a(pp_0_55_0),
    .b(pp_0_55_1),
    .cin(pp_0_55_2),
    .sum(pp_1_55_2),
    .cout(pp_1_56_0)
  );

  MG_FA fa_0_55_1(
    .a(pp_0_55_3),
    .b(pp_0_55_4),
    .cin(pp_0_55_5),
    .sum(pp_1_55_3),
    .cout(pp_1_56_1)
  );

  assign pp_1_56_2 = pp_0_56_0;
  assign pp_1_56_3 = pp_0_56_1;
  assign pp_1_56_4 = pp_0_56_2;
  assign pp_1_56_5 = pp_0_56_3;
  assign pp_1_56_6 = pp_0_56_4;
  assign pp_1_56_7 = pp_0_56_5;
  MG_FA fa_0_57_0(
    .a(pp_0_57_0),
    .b(pp_0_57_1),
    .cin(pp_0_57_2),
    .sum(pp_1_57_0),
    .cout(pp_1_58_0)
  );

  assign pp_1_57_1 = pp_0_57_3;
  assign pp_1_57_2 = pp_0_57_4;
  assign pp_1_58_1 = pp_0_58_0;
  assign pp_1_58_2 = pp_0_58_1;
  assign pp_1_58_3 = pp_0_58_2;
  assign pp_1_58_4 = pp_0_58_3;
  assign pp_1_58_5 = pp_0_58_4;
  MG_FA fa_0_59_0(
    .a(pp_0_59_0),
    .b(pp_0_59_1),
    .cin(pp_0_59_2),
    .sum(pp_1_59_0),
    .cout(pp_1_60_0)
  );

  assign pp_1_59_1 = pp_0_59_3;
  MG_FA fa_0_60_0(
    .a(pp_0_60_0),
    .b(pp_0_60_1),
    .cin(pp_0_60_2),
    .sum(pp_1_60_1),
    .cout(pp_1_61_0)
  );

  assign pp_1_60_2 = pp_0_60_3;
  assign pp_1_61_1 = pp_0_61_0;
  assign pp_1_61_2 = pp_0_61_1;
  assign pp_1_61_3 = pp_0_61_2;
  assign pp_1_62_0 = pp_0_62_0;
  assign pp_1_62_1 = pp_0_62_1;
  assign pp_1_62_2 = pp_0_62_2;
  assign pp_1_63_0 = pp_0_63_0;
  assign pp_1_63_1 = pp_0_63_1;
  assign pp_2_0_0 = pp_1_0_0;
  assign pp_2_0_1 = pp_1_0_1;
  assign pp_2_1_0 = pp_1_1_0;
  assign pp_2_2_0 = pp_1_2_0;
  assign pp_2_2_1 = pp_1_2_1;
  assign pp_2_3_0 = pp_1_3_0;
  assign pp_2_3_1 = pp_1_3_1;
  MG_FA fa_1_4_0(
    .a(pp_1_4_0),
    .b(pp_1_4_1),
    .cin(pp_1_4_2),
    .sum(pp_2_4_0),
    .cout(pp_2_5_0)
  );

  assign pp_2_4_1 = pp_1_4_3;
  assign pp_2_4_2 = pp_1_4_4;
  MG_FA fa_1_5_0(
    .a(pp_1_5_0),
    .b(pp_1_5_1),
    .cin(pp_1_5_2),
    .sum(pp_2_5_1),
    .cout(pp_2_6_0)
  );

  MG_FA fa_1_6_0(
    .a(pp_1_6_0),
    .b(pp_1_6_1),
    .cin(pp_1_6_2),
    .sum(pp_2_6_1),
    .cout(pp_2_7_0)
  );

  MG_FA fa_1_7_0(
    .a(pp_1_7_0),
    .b(pp_1_7_1),
    .cin(pp_1_7_2),
    .sum(pp_2_7_1),
    .cout(pp_2_8_0)
  );

  MG_FA fa_1_8_0(
    .a(pp_1_8_0),
    .b(pp_1_8_1),
    .cin(pp_1_8_2),
    .sum(pp_2_8_1),
    .cout(pp_2_9_0)
  );

  MG_FA fa_1_9_0(
    .a(pp_1_9_0),
    .b(pp_1_9_1),
    .cin(pp_1_9_2),
    .sum(pp_2_9_1),
    .cout(pp_2_10_0)
  );

  MG_FA fa_1_9_1(
    .a(pp_1_9_3),
    .b(pp_1_9_4),
    .cin(pp_1_9_5),
    .sum(pp_2_9_2),
    .cout(pp_2_10_1)
  );

  assign pp_2_9_3 = pp_1_9_6;
  MG_FA fa_1_10_0(
    .a(pp_1_10_0),
    .b(pp_1_10_1),
    .cin(pp_1_10_2),
    .sum(pp_2_10_2),
    .cout(pp_2_11_0)
  );

  MG_FA fa_1_11_0(
    .a(pp_1_11_0),
    .b(pp_1_11_1),
    .cin(pp_1_11_2),
    .sum(pp_2_11_1),
    .cout(pp_2_12_0)
  );

  assign pp_2_11_2 = pp_1_11_3;
  MG_FA fa_1_12_0(
    .a(pp_1_12_0),
    .b(pp_1_12_1),
    .cin(pp_1_12_2),
    .sum(pp_2_12_1),
    .cout(pp_2_13_0)
  );

  MG_FA fa_1_12_1(
    .a(pp_1_12_3),
    .b(pp_1_12_4),
    .cin(pp_1_12_5),
    .sum(pp_2_12_2),
    .cout(pp_2_13_1)
  );

  MG_FA fa_1_13_0(
    .a(pp_1_13_0),
    .b(pp_1_13_1),
    .cin(pp_1_13_2),
    .sum(pp_2_13_2),
    .cout(pp_2_14_0)
  );

  MG_FA fa_1_13_1(
    .a(pp_1_13_3),
    .b(pp_1_13_4),
    .cin(pp_1_13_5),
    .sum(pp_2_13_3),
    .cout(pp_2_14_1)
  );

  assign pp_2_13_4 = pp_1_13_6;
  MG_FA fa_1_14_0(
    .a(pp_1_14_0),
    .b(pp_1_14_1),
    .cin(pp_1_14_2),
    .sum(pp_2_14_2),
    .cout(pp_2_15_0)
  );

  assign pp_2_14_3 = pp_1_14_3;
  MG_FA fa_1_15_0(
    .a(pp_1_15_0),
    .b(pp_1_15_1),
    .cin(pp_1_15_2),
    .sum(pp_2_15_1),
    .cout(pp_2_16_0)
  );

  MG_FA fa_1_15_1(
    .a(pp_1_15_3),
    .b(pp_1_15_4),
    .cin(pp_1_15_5),
    .sum(pp_2_15_2),
    .cout(pp_2_16_1)
  );

  assign pp_2_15_3 = pp_1_15_6;
  MG_FA fa_1_16_0(
    .a(pp_1_16_0),
    .b(pp_1_16_1),
    .cin(pp_1_16_2),
    .sum(pp_2_16_2),
    .cout(pp_2_17_0)
  );

  MG_FA fa_1_16_1(
    .a(pp_1_16_3),
    .b(pp_1_16_4),
    .cin(pp_1_16_5),
    .sum(pp_2_16_3),
    .cout(pp_2_17_1)
  );

  MG_FA fa_1_17_0(
    .a(pp_1_17_0),
    .b(pp_1_17_1),
    .cin(pp_1_17_2),
    .sum(pp_2_17_2),
    .cout(pp_2_18_0)
  );

  MG_FA fa_1_17_1(
    .a(pp_1_17_3),
    .b(pp_1_17_4),
    .cin(pp_1_17_5),
    .sum(pp_2_17_3),
    .cout(pp_2_18_1)
  );

  MG_FA fa_1_18_0(
    .a(pp_1_18_0),
    .b(pp_1_18_1),
    .cin(pp_1_18_2),
    .sum(pp_2_18_2),
    .cout(pp_2_19_0)
  );

  MG_FA fa_1_18_1(
    .a(pp_1_18_3),
    .b(pp_1_18_4),
    .cin(pp_1_18_5),
    .sum(pp_2_18_3),
    .cout(pp_2_19_1)
  );

  MG_FA fa_1_18_2(
    .a(pp_1_18_6),
    .b(pp_1_18_7),
    .cin(pp_1_18_8),
    .sum(pp_2_18_4),
    .cout(pp_2_19_2)
  );

  assign pp_2_18_5 = pp_1_18_9;
  MG_FA fa_1_19_0(
    .a(pp_1_19_0),
    .b(pp_1_19_1),
    .cin(pp_1_19_2),
    .sum(pp_2_19_3),
    .cout(pp_2_20_0)
  );

  MG_FA fa_1_19_1(
    .a(pp_1_19_3),
    .b(pp_1_19_4),
    .cin(pp_1_19_5),
    .sum(pp_2_19_4),
    .cout(pp_2_20_1)
  );

  MG_FA fa_1_20_0(
    .a(pp_1_20_0),
    .b(pp_1_20_1),
    .cin(pp_1_20_2),
    .sum(pp_2_20_2),
    .cout(pp_2_21_0)
  );

  MG_FA fa_1_20_1(
    .a(pp_1_20_3),
    .b(pp_1_20_4),
    .cin(pp_1_20_5),
    .sum(pp_2_20_3),
    .cout(pp_2_21_1)
  );

  assign pp_2_20_4 = pp_1_20_6;
  MG_FA fa_1_21_0(
    .a(pp_1_21_0),
    .b(pp_1_21_1),
    .cin(pp_1_21_2),
    .sum(pp_2_21_2),
    .cout(pp_2_22_0)
  );

  MG_FA fa_1_21_1(
    .a(pp_1_21_3),
    .b(pp_1_21_4),
    .cin(pp_1_21_5),
    .sum(pp_2_21_3),
    .cout(pp_2_22_1)
  );

  MG_FA fa_1_21_2(
    .a(pp_1_21_6),
    .b(pp_1_21_7),
    .cin(pp_1_21_8),
    .sum(pp_2_21_4),
    .cout(pp_2_22_2)
  );

  MG_FA fa_1_22_0(
    .a(pp_1_22_0),
    .b(pp_1_22_1),
    .cin(pp_1_22_2),
    .sum(pp_2_22_3),
    .cout(pp_2_23_0)
  );

  MG_FA fa_1_22_1(
    .a(pp_1_22_3),
    .b(pp_1_22_4),
    .cin(pp_1_22_5),
    .sum(pp_2_22_4),
    .cout(pp_2_23_1)
  );

  MG_HA ha_1_22_2(
    .a(pp_1_22_6),
    .b(pp_1_22_7),
    .sum(pp_2_22_5),
    .cout(pp_2_23_2)
  );

  MG_FA fa_1_23_0(
    .a(pp_1_23_0),
    .b(pp_1_23_1),
    .cin(pp_1_23_2),
    .sum(pp_2_23_3),
    .cout(pp_2_24_0)
  );

  MG_FA fa_1_23_1(
    .a(pp_1_23_3),
    .b(pp_1_23_4),
    .cin(pp_1_23_5),
    .sum(pp_2_23_4),
    .cout(pp_2_24_1)
  );

  assign pp_2_23_5 = pp_1_23_6;
  assign pp_2_23_6 = pp_1_23_7;
  assign pp_2_24_2 = pp_1_24_0;
  assign pp_2_24_3 = pp_1_24_1;
  assign pp_2_24_4 = pp_1_24_2;
  assign pp_2_24_5 = pp_1_24_3;
  assign pp_2_24_6 = pp_1_24_4;
  assign pp_2_24_7 = pp_1_24_5;
  assign pp_2_24_8 = pp_1_24_6;
  assign pp_2_24_9 = pp_1_24_7;
  assign pp_2_24_10 = pp_1_24_8;
  assign pp_2_24_11 = pp_1_24_9;
  MG_FA fa_1_25_0(
    .a(pp_1_25_0),
    .b(pp_1_25_1),
    .cin(pp_1_25_2),
    .sum(pp_2_25_0),
    .cout(pp_2_26_0)
  );

  MG_FA fa_1_25_1(
    .a(pp_1_25_3),
    .b(pp_1_25_4),
    .cin(pp_1_25_5),
    .sum(pp_2_25_1),
    .cout(pp_2_26_1)
  );

  MG_FA fa_1_25_2(
    .a(pp_1_25_6),
    .b(pp_1_25_7),
    .cin(pp_1_25_8),
    .sum(pp_2_25_2),
    .cout(pp_2_26_2)
  );

  MG_FA fa_1_26_0(
    .a(pp_1_26_0),
    .b(pp_1_26_1),
    .cin(pp_1_26_2),
    .sum(pp_2_26_3),
    .cout(pp_2_27_0)
  );

  MG_FA fa_1_26_1(
    .a(pp_1_26_3),
    .b(pp_1_26_4),
    .cin(pp_1_26_5),
    .sum(pp_2_26_4),
    .cout(pp_2_27_1)
  );

  MG_FA fa_1_26_2(
    .a(pp_1_26_6),
    .b(pp_1_26_7),
    .cin(pp_1_26_8),
    .sum(pp_2_26_5),
    .cout(pp_2_27_2)
  );

  MG_FA fa_1_27_0(
    .a(pp_1_27_0),
    .b(pp_1_27_1),
    .cin(pp_1_27_2),
    .sum(pp_2_27_3),
    .cout(pp_2_28_0)
  );

  MG_FA fa_1_27_1(
    .a(pp_1_27_3),
    .b(pp_1_27_4),
    .cin(pp_1_27_5),
    .sum(pp_2_27_4),
    .cout(pp_2_28_1)
  );

  MG_FA fa_1_27_2(
    .a(pp_1_27_6),
    .b(pp_1_27_7),
    .cin(pp_1_27_8),
    .sum(pp_2_27_5),
    .cout(pp_2_28_2)
  );

  MG_FA fa_1_27_3(
    .a(pp_1_27_9),
    .b(pp_1_27_10),
    .cin(pp_1_27_11),
    .sum(pp_2_27_6),
    .cout(pp_2_28_3)
  );

  assign pp_2_27_7 = pp_1_27_12;
  MG_FA fa_1_28_0(
    .a(pp_1_28_0),
    .b(pp_1_28_1),
    .cin(pp_1_28_2),
    .sum(pp_2_28_4),
    .cout(pp_2_29_0)
  );

  MG_FA fa_1_28_1(
    .a(pp_1_28_3),
    .b(pp_1_28_4),
    .cin(pp_1_28_5),
    .sum(pp_2_28_5),
    .cout(pp_2_29_1)
  );

  MG_FA fa_1_28_2(
    .a(pp_1_28_6),
    .b(pp_1_28_7),
    .cin(pp_1_28_8),
    .sum(pp_2_28_6),
    .cout(pp_2_29_2)
  );

  MG_FA fa_1_29_0(
    .a(pp_1_29_0),
    .b(pp_1_29_1),
    .cin(pp_1_29_2),
    .sum(pp_2_29_3),
    .cout(pp_2_30_0)
  );

  MG_FA fa_1_29_1(
    .a(pp_1_29_3),
    .b(pp_1_29_4),
    .cin(pp_1_29_5),
    .sum(pp_2_29_4),
    .cout(pp_2_30_1)
  );

  MG_FA fa_1_29_2(
    .a(pp_1_29_6),
    .b(pp_1_29_7),
    .cin(pp_1_29_8),
    .sum(pp_2_29_5),
    .cout(pp_2_30_2)
  );

  assign pp_2_29_6 = pp_1_29_9;
  MG_FA fa_1_30_0(
    .a(pp_1_30_0),
    .b(pp_1_30_1),
    .cin(pp_1_30_2),
    .sum(pp_2_30_3),
    .cout(pp_2_31_0)
  );

  MG_FA fa_1_30_1(
    .a(pp_1_30_3),
    .b(pp_1_30_4),
    .cin(pp_1_30_5),
    .sum(pp_2_30_4),
    .cout(pp_2_31_1)
  );

  MG_FA fa_1_30_2(
    .a(pp_1_30_6),
    .b(pp_1_30_7),
    .cin(pp_1_30_8),
    .sum(pp_2_30_5),
    .cout(pp_2_31_2)
  );

  MG_FA fa_1_30_3(
    .a(pp_1_30_9),
    .b(pp_1_30_10),
    .cin(pp_1_30_11),
    .sum(pp_2_30_6),
    .cout(pp_2_31_3)
  );

  MG_FA fa_1_31_0(
    .a(pp_1_31_0),
    .b(pp_1_31_1),
    .cin(pp_1_31_2),
    .sum(pp_2_31_4),
    .cout(pp_2_32_0)
  );

  MG_FA fa_1_31_1(
    .a(pp_1_31_3),
    .b(pp_1_31_4),
    .cin(pp_1_31_5),
    .sum(pp_2_31_5),
    .cout(pp_2_32_1)
  );

  MG_FA fa_1_31_2(
    .a(pp_1_31_6),
    .b(pp_1_31_7),
    .cin(pp_1_31_8),
    .sum(pp_2_31_6),
    .cout(pp_2_32_2)
  );

  MG_FA fa_1_31_3(
    .a(pp_1_31_9),
    .b(pp_1_31_10),
    .cin(pp_1_31_11),
    .sum(pp_2_31_7),
    .cout(pp_2_32_3)
  );

  MG_FA fa_1_32_0(
    .a(pp_1_32_0),
    .b(pp_1_32_1),
    .cin(pp_1_32_2),
    .sum(pp_2_32_4),
    .cout(pp_2_33_0)
  );

  MG_FA fa_1_32_1(
    .a(pp_1_32_3),
    .b(pp_1_32_4),
    .cin(pp_1_32_5),
    .sum(pp_2_32_5),
    .cout(pp_2_33_1)
  );

  assign pp_2_32_6 = pp_1_32_6;
  assign pp_2_32_7 = pp_1_32_7;
  assign pp_2_32_8 = pp_1_32_8;
  assign pp_2_32_9 = pp_1_32_9;
  assign pp_2_32_10 = pp_1_32_10;
  assign pp_2_32_11 = pp_1_32_11;
  MG_FA fa_1_33_0(
    .a(pp_1_33_0),
    .b(pp_1_33_1),
    .cin(pp_1_33_2),
    .sum(pp_2_33_2),
    .cout(pp_2_34_0)
  );

  MG_FA fa_1_33_1(
    .a(pp_1_33_3),
    .b(pp_1_33_4),
    .cin(pp_1_33_5),
    .sum(pp_2_33_3),
    .cout(pp_2_34_1)
  );

  MG_FA fa_1_33_2(
    .a(pp_1_33_10),
    .b(pp_1_33_11),
    .cin(pp_1_33_8),
    .sum(pp_2_33_4),
    .cout(pp_2_34_2)
  );

  MG_FA fa_1_33_3(
    .a(pp_1_33_9),
    .b(pp_1_33_6),
    .cin(pp_1_33_7),
    .sum(pp_2_33_5),
    .cout(pp_2_34_3)
  );

  MG_FA fa_1_34_0(
    .a(pp_1_34_0),
    .b(pp_1_34_1),
    .cin(pp_1_34_2),
    .sum(pp_2_34_4),
    .cout(pp_2_35_0)
  );

  MG_FA fa_1_34_1(
    .a(pp_1_34_3),
    .b(pp_1_34_4),
    .cin(pp_1_34_5),
    .sum(pp_2_34_5),
    .cout(pp_2_35_1)
  );

  MG_FA fa_1_34_2(
    .a(pp_1_34_6),
    .b(pp_1_34_7),
    .cin(pp_1_34_8),
    .sum(pp_2_34_6),
    .cout(pp_2_35_2)
  );

  MG_FA fa_1_34_3(
    .a(pp_1_34_9),
    .b(pp_1_34_10),
    .cin(pp_1_34_11),
    .sum(pp_2_34_7),
    .cout(pp_2_35_3)
  );

  MG_FA fa_1_35_0(
    .a(pp_1_35_0),
    .b(pp_1_35_1),
    .cin(pp_1_35_2),
    .sum(pp_2_35_4),
    .cout(pp_2_36_0)
  );

  MG_FA fa_1_35_1(
    .a(pp_1_35_3),
    .b(pp_1_35_4),
    .cin(pp_1_35_5),
    .sum(pp_2_35_5),
    .cout(pp_2_36_1)
  );

  MG_FA fa_1_35_2(
    .a(pp_1_35_6),
    .b(pp_1_35_7),
    .cin(pp_1_35_8),
    .sum(pp_2_35_6),
    .cout(pp_2_36_2)
  );

  MG_FA fa_1_35_3(
    .a(pp_1_35_9),
    .b(pp_1_35_10),
    .cin(pp_1_35_11),
    .sum(pp_2_35_7),
    .cout(pp_2_36_3)
  );

  MG_FA fa_1_36_0(
    .a(pp_1_36_0),
    .b(pp_1_36_1),
    .cin(pp_1_36_2),
    .sum(pp_2_36_4),
    .cout(pp_2_37_0)
  );

  MG_FA fa_1_36_1(
    .a(pp_1_36_3),
    .b(pp_1_36_4),
    .cin(pp_1_36_5),
    .sum(pp_2_36_5),
    .cout(pp_2_37_1)
  );

  MG_FA fa_1_36_2(
    .a(pp_1_36_6),
    .b(pp_1_36_7),
    .cin(pp_1_36_8),
    .sum(pp_2_36_6),
    .cout(pp_2_37_2)
  );

  assign pp_2_36_7 = pp_1_36_9;
  assign pp_2_36_8 = pp_1_36_10;
  MG_FA fa_1_37_0(
    .a(pp_1_37_0),
    .b(pp_1_37_1),
    .cin(pp_1_37_2),
    .sum(pp_2_37_3),
    .cout(pp_2_38_0)
  );

  MG_FA fa_1_37_1(
    .a(pp_1_37_3),
    .b(pp_1_37_4),
    .cin(pp_1_37_5),
    .sum(pp_2_37_4),
    .cout(pp_2_38_1)
  );

  MG_FA fa_1_37_2(
    .a(pp_1_37_6),
    .b(pp_1_37_7),
    .cin(pp_1_37_8),
    .sum(pp_2_37_5),
    .cout(pp_2_38_2)
  );

  MG_FA fa_1_37_3(
    .a(pp_1_37_9),
    .b(pp_1_37_10),
    .cin(pp_1_37_11),
    .sum(pp_2_37_6),
    .cout(pp_2_38_3)
  );

  MG_FA fa_1_38_0(
    .a(pp_1_38_0),
    .b(pp_1_38_1),
    .cin(pp_1_38_2),
    .sum(pp_2_38_4),
    .cout(pp_2_39_0)
  );

  MG_FA fa_1_38_1(
    .a(pp_1_38_3),
    .b(pp_1_38_4),
    .cin(pp_1_38_5),
    .sum(pp_2_38_5),
    .cout(pp_2_39_1)
  );

  MG_FA fa_1_38_2(
    .a(pp_1_38_6),
    .b(pp_1_38_7),
    .cin(pp_1_38_8),
    .sum(pp_2_38_6),
    .cout(pp_2_39_2)
  );

  MG_FA fa_1_39_0(
    .a(pp_1_39_0),
    .b(pp_1_39_1),
    .cin(pp_1_39_2),
    .sum(pp_2_39_3),
    .cout(pp_2_40_0)
  );

  MG_FA fa_1_39_1(
    .a(pp_1_39_3),
    .b(pp_1_39_4),
    .cin(pp_1_39_5),
    .sum(pp_2_39_4),
    .cout(pp_2_40_1)
  );

  MG_FA fa_1_39_2(
    .a(pp_1_39_6),
    .b(pp_1_39_7),
    .cin(pp_1_39_8),
    .sum(pp_2_39_5),
    .cout(pp_2_40_2)
  );

  assign pp_2_39_6 = pp_1_39_9;
  assign pp_2_39_7 = pp_1_39_10;
  MG_FA fa_1_40_0(
    .a(pp_1_40_0),
    .b(pp_1_40_1),
    .cin(pp_1_40_2),
    .sum(pp_2_40_3),
    .cout(pp_2_41_0)
  );

  MG_FA fa_1_40_1(
    .a(pp_1_40_3),
    .b(pp_1_40_4),
    .cin(pp_1_40_5),
    .sum(pp_2_40_4),
    .cout(pp_2_41_1)
  );

  assign pp_2_40_5 = pp_1_40_6;
  assign pp_2_40_6 = pp_1_40_7;
  assign pp_2_40_7 = pp_1_40_8;
  assign pp_2_40_8 = pp_1_40_9;
  MG_FA fa_1_41_0(
    .a(pp_1_41_0),
    .b(pp_1_41_1),
    .cin(pp_1_41_2),
    .sum(pp_2_41_2),
    .cout(pp_2_42_0)
  );

  MG_FA fa_1_41_1(
    .a(pp_1_41_3),
    .b(pp_1_41_4),
    .cin(pp_1_41_5),
    .sum(pp_2_41_3),
    .cout(pp_2_42_1)
  );

  MG_FA fa_1_41_2(
    .a(pp_1_41_6),
    .b(pp_1_41_7),
    .cin(pp_1_41_8),
    .sum(pp_2_41_4),
    .cout(pp_2_42_2)
  );

  MG_FA fa_1_42_0(
    .a(pp_1_42_0),
    .b(pp_1_42_1),
    .cin(pp_1_42_2),
    .sum(pp_2_42_3),
    .cout(pp_2_43_0)
  );

  MG_FA fa_1_42_1(
    .a(pp_1_42_3),
    .b(pp_1_42_4),
    .cin(pp_1_42_5),
    .sum(pp_2_42_4),
    .cout(pp_2_43_1)
  );

  MG_FA fa_1_42_2(
    .a(pp_1_42_6),
    .b(pp_1_42_7),
    .cin(pp_1_42_8),
    .sum(pp_2_42_5),
    .cout(pp_2_43_2)
  );

  MG_FA fa_1_43_0(
    .a(pp_1_43_0),
    .b(pp_1_43_1),
    .cin(pp_1_43_2),
    .sum(pp_2_43_3),
    .cout(pp_2_44_0)
  );

  MG_FA fa_1_43_1(
    .a(pp_1_43_3),
    .b(pp_1_43_4),
    .cin(pp_1_43_5),
    .sum(pp_2_43_4),
    .cout(pp_2_44_1)
  );

  MG_FA fa_1_43_2(
    .a(pp_1_43_6),
    .b(pp_1_43_7),
    .cin(pp_1_43_8),
    .sum(pp_2_43_5),
    .cout(pp_2_44_2)
  );

  MG_FA fa_1_43_3(
    .a(pp_1_43_9),
    .b(pp_1_43_10),
    .cin(pp_1_43_11),
    .sum(pp_2_43_6),
    .cout(pp_2_44_3)
  );

  MG_FA fa_1_44_0(
    .a(pp_1_44_0),
    .b(pp_1_44_1),
    .cin(pp_1_44_2),
    .sum(pp_2_44_4),
    .cout(pp_2_45_0)
  );

  MG_FA fa_1_44_1(
    .a(pp_1_44_3),
    .b(pp_1_44_4),
    .cin(pp_1_44_5),
    .sum(pp_2_44_5),
    .cout(pp_2_45_1)
  );

  MG_FA fa_1_45_0(
    .a(pp_1_45_0),
    .b(pp_1_45_1),
    .cin(pp_1_45_2),
    .sum(pp_2_45_2),
    .cout(pp_2_46_0)
  );

  MG_FA fa_1_45_1(
    .a(pp_1_45_3),
    .b(pp_1_45_4),
    .cin(pp_1_45_5),
    .sum(pp_2_45_3),
    .cout(pp_2_46_1)
  );

  MG_FA fa_1_45_2(
    .a(pp_1_45_6),
    .b(pp_1_45_7),
    .cin(pp_1_45_8),
    .sum(pp_2_45_4),
    .cout(pp_2_46_2)
  );

  MG_FA fa_1_45_3(
    .a(pp_1_45_9),
    .b(pp_1_45_10),
    .cin(pp_1_45_11),
    .sum(pp_2_45_5),
    .cout(pp_2_46_3)
  );

  assign pp_2_45_6 = pp_1_45_12;
  MG_FA fa_1_46_0(
    .a(pp_1_46_0),
    .b(pp_1_46_1),
    .cin(pp_1_46_2),
    .sum(pp_2_46_4),
    .cout(pp_2_47_0)
  );

  MG_FA fa_1_46_1(
    .a(pp_1_46_3),
    .b(pp_1_46_4),
    .cin(pp_1_46_5),
    .sum(pp_2_46_5),
    .cout(pp_2_47_1)
  );

  MG_FA fa_1_46_2(
    .a(pp_1_46_6),
    .b(pp_1_46_7),
    .cin(pp_1_46_8),
    .sum(pp_2_46_6),
    .cout(pp_2_47_2)
  );

  MG_FA fa_1_47_0(
    .a(pp_1_47_0),
    .b(pp_1_47_1),
    .cin(pp_1_47_2),
    .sum(pp_2_47_3),
    .cout(pp_2_48_0)
  );

  MG_FA fa_1_47_1(
    .a(pp_1_47_3),
    .b(pp_1_47_4),
    .cin(pp_1_47_5),
    .sum(pp_2_47_4),
    .cout(pp_2_48_1)
  );

  MG_FA fa_1_48_0(
    .a(pp_1_48_0),
    .b(pp_1_48_1),
    .cin(pp_1_48_2),
    .sum(pp_2_48_2),
    .cout(pp_2_49_0)
  );

  MG_FA fa_1_48_1(
    .a(pp_1_48_3),
    .b(pp_1_48_4),
    .cin(pp_1_48_5),
    .sum(pp_2_48_3),
    .cout(pp_2_49_1)
  );

  MG_FA fa_1_48_2(
    .a(pp_1_48_6),
    .b(pp_1_48_7),
    .cin(pp_1_48_8),
    .sum(pp_2_48_4),
    .cout(pp_2_49_2)
  );

  MG_FA fa_1_49_0(
    .a(pp_1_49_0),
    .b(pp_1_49_1),
    .cin(pp_1_49_2),
    .sum(pp_2_49_3),
    .cout(pp_2_50_0)
  );

  assign pp_2_49_4 = pp_1_49_3;
  assign pp_2_49_5 = pp_1_49_4;
  MG_FA fa_1_50_0(
    .a(pp_1_50_0),
    .b(pp_1_50_1),
    .cin(pp_1_50_2),
    .sum(pp_2_50_1),
    .cout(pp_2_51_0)
  );

  MG_FA fa_1_50_1(
    .a(pp_1_50_3),
    .b(pp_1_50_4),
    .cin(pp_1_50_5),
    .sum(pp_2_50_2),
    .cout(pp_2_51_1)
  );

  MG_FA fa_1_51_0(
    .a(pp_1_51_0),
    .b(pp_1_51_1),
    .cin(pp_1_51_2),
    .sum(pp_2_51_2),
    .cout(pp_2_52_0)
  );

  MG_FA fa_1_51_1(
    .a(pp_1_51_3),
    .b(pp_1_51_4),
    .cin(pp_1_51_5),
    .sum(pp_2_51_3),
    .cout(pp_2_52_1)
  );

  assign pp_2_51_4 = pp_1_51_6;
  MG_FA fa_1_52_0(
    .a(pp_1_52_0),
    .b(pp_1_52_1),
    .cin(pp_1_52_2),
    .sum(pp_2_52_2),
    .cout(pp_2_53_0)
  );

  MG_FA fa_1_52_1(
    .a(pp_1_52_3),
    .b(pp_1_52_4),
    .cin(pp_1_52_5),
    .sum(pp_2_52_3),
    .cout(pp_2_53_1)
  );

  MG_FA fa_1_53_0(
    .a(pp_1_53_0),
    .b(pp_1_53_1),
    .cin(pp_1_53_2),
    .sum(pp_2_53_2),
    .cout(pp_2_54_0)
  );

  MG_FA fa_1_53_1(
    .a(pp_1_53_3),
    .b(pp_1_53_4),
    .cin(pp_1_53_5),
    .sum(pp_2_53_3),
    .cout(pp_2_54_1)
  );

  MG_FA fa_1_53_2(
    .a(pp_1_53_6),
    .b(pp_1_53_7),
    .cin(pp_1_53_8),
    .sum(pp_2_53_4),
    .cout(pp_2_54_2)
  );

  MG_FA fa_1_54_0(
    .a(pp_1_54_0),
    .b(pp_1_54_1),
    .cin(pp_1_54_2),
    .sum(pp_2_54_3),
    .cout(pp_2_55_0)
  );

  assign pp_2_55_1 = pp_1_55_0;
  assign pp_2_55_2 = pp_1_55_1;
  assign pp_2_55_3 = pp_1_55_2;
  assign pp_2_55_4 = pp_1_55_3;
  MG_FA fa_1_56_0(
    .a(pp_1_56_0),
    .b(pp_1_56_1),
    .cin(pp_1_56_2),
    .sum(pp_2_56_0),
    .cout(pp_2_57_0)
  );

  assign pp_2_56_1 = pp_1_56_3;
  assign pp_2_56_2 = pp_1_56_4;
  assign pp_2_56_3 = pp_1_56_5;
  assign pp_2_56_4 = pp_1_56_6;
  assign pp_2_56_5 = pp_1_56_7;
  MG_FA fa_1_57_0(
    .a(pp_1_57_0),
    .b(pp_1_57_1),
    .cin(pp_1_57_2),
    .sum(pp_2_57_1),
    .cout(pp_2_58_0)
  );

  MG_FA fa_1_58_0(
    .a(pp_1_58_0),
    .b(pp_1_58_1),
    .cin(pp_1_58_2),
    .sum(pp_2_58_1),
    .cout(pp_2_59_0)
  );

  MG_FA fa_1_58_1(
    .a(pp_1_58_3),
    .b(pp_1_58_4),
    .cin(pp_1_58_5),
    .sum(pp_2_58_2),
    .cout(pp_2_59_1)
  );

  assign pp_2_59_2 = pp_1_59_0;
  assign pp_2_59_3 = pp_1_59_1;
  MG_FA fa_1_60_0(
    .a(pp_1_60_0),
    .b(pp_1_60_1),
    .cin(pp_1_60_2),
    .sum(pp_2_60_0),
    .cout(pp_2_61_0)
  );

  MG_FA fa_1_61_0(
    .a(pp_1_61_0),
    .b(pp_1_61_1),
    .cin(pp_1_61_2),
    .sum(pp_2_61_1),
    .cout(pp_2_62_0)
  );

  assign pp_2_61_2 = pp_1_61_3;
  MG_FA fa_1_62_0(
    .a(pp_1_62_0),
    .b(pp_1_62_1),
    .cin(pp_1_62_2),
    .sum(pp_2_62_1),
    .cout(pp_2_63_0)
  );

  assign pp_2_63_1 = pp_1_63_0;
  assign pp_2_63_2 = pp_1_63_1;
  assign pp_3_0_0 = pp_2_0_0;
  assign pp_3_0_1 = pp_2_0_1;
  assign pp_3_1_0 = pp_2_1_0;
  assign pp_3_2_0 = pp_2_2_0;
  assign pp_3_2_1 = pp_2_2_1;
  assign pp_3_3_0 = pp_2_3_0;
  assign pp_3_3_1 = pp_2_3_1;
  assign pp_3_4_0 = pp_2_4_0;
  assign pp_3_4_1 = pp_2_4_1;
  assign pp_3_4_2 = pp_2_4_2;
  MG_HA ha_2_5_0(
    .a(pp_2_5_0),
    .b(pp_2_5_1),
    .sum(pp_3_5_0),
    .cout(pp_3_6_0)
  );

  assign pp_3_6_1 = pp_2_6_0;
  assign pp_3_6_2 = pp_2_6_1;
  MG_HA ha_2_7_0(
    .a(pp_2_7_0),
    .b(pp_2_7_1),
    .sum(pp_3_7_0),
    .cout(pp_3_8_0)
  );

  assign pp_3_8_1 = pp_2_8_0;
  assign pp_3_8_2 = pp_2_8_1;
  assign pp_3_9_0 = pp_2_9_0;
  assign pp_3_9_1 = pp_2_9_1;
  assign pp_3_9_2 = pp_2_9_2;
  assign pp_3_9_3 = pp_2_9_3;
  MG_FA fa_2_10_0(
    .a(pp_2_10_0),
    .b(pp_2_10_1),
    .cin(pp_2_10_2),
    .sum(pp_3_10_0),
    .cout(pp_3_11_0)
  );

  MG_FA fa_2_11_0(
    .a(pp_2_11_0),
    .b(pp_2_11_1),
    .cin(pp_2_11_2),
    .sum(pp_3_11_1),
    .cout(pp_3_12_0)
  );

  MG_FA fa_2_12_0(
    .a(pp_2_12_0),
    .b(pp_2_12_1),
    .cin(pp_2_12_2),
    .sum(pp_3_12_1),
    .cout(pp_3_13_0)
  );

  MG_FA fa_2_13_0(
    .a(pp_2_13_0),
    .b(pp_2_13_1),
    .cin(pp_2_13_2),
    .sum(pp_3_13_1),
    .cout(pp_3_14_0)
  );

  assign pp_3_13_2 = pp_2_13_3;
  assign pp_3_13_3 = pp_2_13_4;
  MG_FA fa_2_14_0(
    .a(pp_2_14_0),
    .b(pp_2_14_1),
    .cin(pp_2_14_2),
    .sum(pp_3_14_1),
    .cout(pp_3_15_0)
  );

  assign pp_3_14_2 = pp_2_14_3;
  MG_FA fa_2_15_0(
    .a(pp_2_15_0),
    .b(pp_2_15_1),
    .cin(pp_2_15_2),
    .sum(pp_3_15_1),
    .cout(pp_3_16_0)
  );

  assign pp_3_15_2 = pp_2_15_3;
  MG_HA ha_2_16_0(
    .a(pp_2_16_0),
    .b(pp_2_16_1),
    .sum(pp_3_16_1),
    .cout(pp_3_17_0)
  );

  assign pp_3_16_2 = pp_2_16_2;
  assign pp_3_16_3 = pp_2_16_3;
  MG_FA fa_2_17_0(
    .a(pp_2_17_0),
    .b(pp_2_17_1),
    .cin(pp_2_17_2),
    .sum(pp_3_17_1),
    .cout(pp_3_18_0)
  );

  assign pp_3_17_2 = pp_2_17_3;
  MG_FA fa_2_18_0(
    .a(pp_2_18_0),
    .b(pp_2_18_1),
    .cin(pp_2_18_2),
    .sum(pp_3_18_1),
    .cout(pp_3_19_0)
  );

  MG_FA fa_2_18_1(
    .a(pp_2_18_3),
    .b(pp_2_18_4),
    .cin(pp_2_18_5),
    .sum(pp_3_18_2),
    .cout(pp_3_19_1)
  );

  MG_FA fa_2_19_0(
    .a(pp_2_19_0),
    .b(pp_2_19_1),
    .cin(pp_2_19_2),
    .sum(pp_3_19_2),
    .cout(pp_3_20_0)
  );

  MG_HA ha_2_19_1(
    .a(pp_2_19_3),
    .b(pp_2_19_4),
    .sum(pp_3_19_3),
    .cout(pp_3_20_1)
  );

  MG_FA fa_2_20_0(
    .a(pp_2_20_0),
    .b(pp_2_20_1),
    .cin(pp_2_20_2),
    .sum(pp_3_20_2),
    .cout(pp_3_21_0)
  );

  MG_HA ha_2_20_1(
    .a(pp_2_20_3),
    .b(pp_2_20_4),
    .sum(pp_3_20_3),
    .cout(pp_3_21_1)
  );

  MG_FA fa_2_21_0(
    .a(pp_2_21_0),
    .b(pp_2_21_1),
    .cin(pp_2_21_2),
    .sum(pp_3_21_2),
    .cout(pp_3_22_0)
  );

  MG_HA ha_2_21_1(
    .a(pp_2_21_3),
    .b(pp_2_21_4),
    .sum(pp_3_21_3),
    .cout(pp_3_22_1)
  );

  MG_FA fa_2_22_0(
    .a(pp_2_22_0),
    .b(pp_2_22_1),
    .cin(pp_2_22_2),
    .sum(pp_3_22_2),
    .cout(pp_3_23_0)
  );

  assign pp_3_22_3 = pp_2_22_3;
  assign pp_3_22_4 = pp_2_22_4;
  assign pp_3_22_5 = pp_2_22_5;
  MG_FA fa_2_23_0(
    .a(pp_2_23_0),
    .b(pp_2_23_1),
    .cin(pp_2_23_2),
    .sum(pp_3_23_1),
    .cout(pp_3_24_0)
  );

  MG_FA fa_2_23_1(
    .a(pp_2_23_3),
    .b(pp_2_23_4),
    .cin(pp_2_23_5),
    .sum(pp_3_23_2),
    .cout(pp_3_24_1)
  );

  assign pp_3_23_3 = pp_2_23_6;
  MG_FA fa_2_24_0(
    .a(pp_2_24_0),
    .b(pp_2_24_1),
    .cin(pp_2_24_2),
    .sum(pp_3_24_2),
    .cout(pp_3_25_0)
  );

  MG_FA fa_2_24_1(
    .a(pp_2_24_3),
    .b(pp_2_24_4),
    .cin(pp_2_24_5),
    .sum(pp_3_24_3),
    .cout(pp_3_25_1)
  );

  MG_FA fa_2_24_2(
    .a(pp_2_24_6),
    .b(pp_2_24_7),
    .cin(pp_2_24_8),
    .sum(pp_3_24_4),
    .cout(pp_3_25_2)
  );

  MG_FA fa_2_24_3(
    .a(pp_2_24_9),
    .b(pp_2_24_10),
    .cin(pp_2_24_11),
    .sum(pp_3_24_5),
    .cout(pp_3_25_3)
  );

  MG_HA ha_2_25_0(
    .a(pp_2_25_0),
    .b(pp_2_25_1),
    .sum(pp_3_25_4),
    .cout(pp_3_26_0)
  );

  assign pp_3_25_5 = pp_2_25_2;
  MG_FA fa_2_26_0(
    .a(pp_2_26_0),
    .b(pp_2_26_1),
    .cin(pp_2_26_2),
    .sum(pp_3_26_1),
    .cout(pp_3_27_0)
  );

  MG_FA fa_2_26_1(
    .a(pp_2_26_3),
    .b(pp_2_26_4),
    .cin(pp_2_26_5),
    .sum(pp_3_26_2),
    .cout(pp_3_27_1)
  );

  MG_FA fa_2_27_0(
    .a(pp_2_27_0),
    .b(pp_2_27_1),
    .cin(pp_2_27_2),
    .sum(pp_3_27_2),
    .cout(pp_3_28_0)
  );

  MG_FA fa_2_27_1(
    .a(pp_2_27_3),
    .b(pp_2_27_4),
    .cin(pp_2_27_5),
    .sum(pp_3_27_3),
    .cout(pp_3_28_1)
  );

  assign pp_3_27_4 = pp_2_27_6;
  assign pp_3_27_5 = pp_2_27_7;
  MG_FA fa_2_28_0(
    .a(pp_2_28_0),
    .b(pp_2_28_1),
    .cin(pp_2_28_2),
    .sum(pp_3_28_2),
    .cout(pp_3_29_0)
  );

  MG_FA fa_2_28_1(
    .a(pp_2_28_3),
    .b(pp_2_28_4),
    .cin(pp_2_28_5),
    .sum(pp_3_28_3),
    .cout(pp_3_29_1)
  );

  assign pp_3_28_4 = pp_2_28_6;
  MG_FA fa_2_29_0(
    .a(pp_2_29_0),
    .b(pp_2_29_1),
    .cin(pp_2_29_2),
    .sum(pp_3_29_2),
    .cout(pp_3_30_0)
  );

  MG_FA fa_2_29_1(
    .a(pp_2_29_3),
    .b(pp_2_29_4),
    .cin(pp_2_29_5),
    .sum(pp_3_29_3),
    .cout(pp_3_30_1)
  );

  assign pp_3_29_4 = pp_2_29_6;
  MG_FA fa_2_30_0(
    .a(pp_2_30_0),
    .b(pp_2_30_1),
    .cin(pp_2_30_2),
    .sum(pp_3_30_2),
    .cout(pp_3_31_0)
  );

  MG_HA ha_2_30_1(
    .a(pp_2_30_3),
    .b(pp_2_30_4),
    .sum(pp_3_30_3),
    .cout(pp_3_31_1)
  );

  assign pp_3_30_4 = pp_2_30_5;
  assign pp_3_30_5 = pp_2_30_6;
  MG_FA fa_2_31_0(
    .a(pp_2_31_0),
    .b(pp_2_31_1),
    .cin(pp_2_31_2),
    .sum(pp_3_31_2),
    .cout(pp_3_32_0)
  );

  MG_FA fa_2_31_1(
    .a(pp_2_31_3),
    .b(pp_2_31_4),
    .cin(pp_2_31_5),
    .sum(pp_3_31_3),
    .cout(pp_3_32_1)
  );

  assign pp_3_31_4 = pp_2_31_6;
  assign pp_3_31_5 = pp_2_31_7;
  MG_FA fa_2_32_0(
    .a(pp_2_32_0),
    .b(pp_2_32_1),
    .cin(pp_2_32_2),
    .sum(pp_3_32_2),
    .cout(pp_3_33_0)
  );

  MG_FA fa_2_32_1(
    .a(pp_2_32_3),
    .b(pp_2_32_4),
    .cin(pp_2_32_5),
    .sum(pp_3_32_3),
    .cout(pp_3_33_1)
  );

  MG_FA fa_2_32_2(
    .a(pp_2_32_6),
    .b(pp_2_32_7),
    .cin(pp_2_32_8),
    .sum(pp_3_32_4),
    .cout(pp_3_33_2)
  );

  MG_FA fa_2_32_3(
    .a(pp_2_32_9),
    .b(pp_2_32_10),
    .cin(pp_2_32_11),
    .sum(pp_3_32_5),
    .cout(pp_3_33_3)
  );

  MG_FA fa_2_33_0(
    .a(pp_2_33_0),
    .b(pp_2_33_1),
    .cin(pp_2_33_2),
    .sum(pp_3_33_4),
    .cout(pp_3_34_0)
  );

  MG_FA fa_2_33_1(
    .a(pp_2_33_3),
    .b(pp_2_33_4),
    .cin(pp_2_33_5),
    .sum(pp_3_33_5),
    .cout(pp_3_34_1)
  );

  MG_FA fa_2_34_0(
    .a(pp_2_34_0),
    .b(pp_2_34_1),
    .cin(pp_2_34_2),
    .sum(pp_3_34_2),
    .cout(pp_3_35_0)
  );

  MG_FA fa_2_34_1(
    .a(pp_2_34_3),
    .b(pp_2_34_4),
    .cin(pp_2_34_5),
    .sum(pp_3_34_3),
    .cout(pp_3_35_1)
  );

  assign pp_3_34_4 = pp_2_34_6;
  assign pp_3_34_5 = pp_2_34_7;
  MG_FA fa_2_35_0(
    .a(pp_2_35_0),
    .b(pp_2_35_1),
    .cin(pp_2_35_2),
    .sum(pp_3_35_2),
    .cout(pp_3_36_0)
  );

  MG_FA fa_2_35_1(
    .a(pp_2_35_3),
    .b(pp_2_35_4),
    .cin(pp_2_35_5),
    .sum(pp_3_35_3),
    .cout(pp_3_36_1)
  );

  assign pp_3_35_4 = pp_2_35_6;
  assign pp_3_35_5 = pp_2_35_7;
  MG_FA fa_2_36_0(
    .a(pp_2_36_0),
    .b(pp_2_36_1),
    .cin(pp_2_36_2),
    .sum(pp_3_36_2),
    .cout(pp_3_37_0)
  );

  MG_FA fa_2_36_1(
    .a(pp_2_36_3),
    .b(pp_2_36_4),
    .cin(pp_2_36_5),
    .sum(pp_3_36_3),
    .cout(pp_3_37_1)
  );

  MG_FA fa_2_36_2(
    .a(pp_2_36_6),
    .b(pp_2_36_7),
    .cin(pp_2_36_8),
    .sum(pp_3_36_4),
    .cout(pp_3_37_2)
  );

  MG_FA fa_2_37_0(
    .a(pp_2_37_0),
    .b(pp_2_37_1),
    .cin(pp_2_37_2),
    .sum(pp_3_37_3),
    .cout(pp_3_38_0)
  );

  MG_FA fa_2_37_1(
    .a(pp_2_37_3),
    .b(pp_2_37_4),
    .cin(pp_2_37_5),
    .sum(pp_3_37_4),
    .cout(pp_3_38_1)
  );

  assign pp_3_37_5 = pp_2_37_6;
  MG_FA fa_2_38_0(
    .a(pp_2_38_0),
    .b(pp_2_38_1),
    .cin(pp_2_38_2),
    .sum(pp_3_38_2),
    .cout(pp_3_39_0)
  );

  MG_HA ha_2_38_1(
    .a(pp_2_38_3),
    .b(pp_2_38_4),
    .sum(pp_3_38_3),
    .cout(pp_3_39_1)
  );

  assign pp_3_38_4 = pp_2_38_5;
  assign pp_3_38_5 = pp_2_38_6;
  MG_FA fa_2_39_0(
    .a(pp_2_39_0),
    .b(pp_2_39_1),
    .cin(pp_2_39_2),
    .sum(pp_3_39_2),
    .cout(pp_3_40_0)
  );

  MG_FA fa_2_39_1(
    .a(pp_2_39_3),
    .b(pp_2_39_4),
    .cin(pp_2_39_5),
    .sum(pp_3_39_3),
    .cout(pp_3_40_1)
  );

  assign pp_3_39_4 = pp_2_39_6;
  assign pp_3_39_5 = pp_2_39_7;
  MG_FA fa_2_40_0(
    .a(pp_2_40_0),
    .b(pp_2_40_1),
    .cin(pp_2_40_2),
    .sum(pp_3_40_2),
    .cout(pp_3_41_0)
  );

  MG_FA fa_2_40_1(
    .a(pp_2_40_3),
    .b(pp_2_40_4),
    .cin(pp_2_40_5),
    .sum(pp_3_40_3),
    .cout(pp_3_41_1)
  );

  MG_FA fa_2_40_2(
    .a(pp_2_40_6),
    .b(pp_2_40_7),
    .cin(pp_2_40_8),
    .sum(pp_3_40_4),
    .cout(pp_3_41_2)
  );

  MG_FA fa_2_41_0(
    .a(pp_2_41_0),
    .b(pp_2_41_1),
    .cin(pp_2_41_2),
    .sum(pp_3_41_3),
    .cout(pp_3_42_0)
  );

  assign pp_3_41_4 = pp_2_41_3;
  assign pp_3_41_5 = pp_2_41_4;
  MG_FA fa_2_42_0(
    .a(pp_2_42_0),
    .b(pp_2_42_1),
    .cin(pp_2_42_2),
    .sum(pp_3_42_1),
    .cout(pp_3_43_0)
  );

  MG_FA fa_2_42_1(
    .a(pp_2_42_3),
    .b(pp_2_42_4),
    .cin(pp_2_42_5),
    .sum(pp_3_42_2),
    .cout(pp_3_43_1)
  );

  MG_FA fa_2_43_0(
    .a(pp_2_43_0),
    .b(pp_2_43_1),
    .cin(pp_2_43_2),
    .sum(pp_3_43_2),
    .cout(pp_3_44_0)
  );

  MG_FA fa_2_43_1(
    .a(pp_2_43_3),
    .b(pp_2_43_4),
    .cin(pp_2_43_5),
    .sum(pp_3_43_3),
    .cout(pp_3_44_1)
  );

  assign pp_3_43_4 = pp_2_43_6;
  MG_FA fa_2_44_0(
    .a(pp_2_44_0),
    .b(pp_2_44_1),
    .cin(pp_2_44_2),
    .sum(pp_3_44_2),
    .cout(pp_3_45_0)
  );

  assign pp_3_44_3 = pp_2_44_3;
  assign pp_3_44_4 = pp_2_44_4;
  assign pp_3_44_5 = pp_2_44_5;
  MG_FA fa_2_45_0(
    .a(pp_2_45_0),
    .b(pp_2_45_1),
    .cin(pp_2_45_2),
    .sum(pp_3_45_1),
    .cout(pp_3_46_0)
  );

  MG_FA fa_2_45_1(
    .a(pp_2_45_3),
    .b(pp_2_45_4),
    .cin(pp_2_45_5),
    .sum(pp_3_45_2),
    .cout(pp_3_46_1)
  );

  assign pp_3_45_3 = pp_2_45_6;
  assign pp_3_46_2 = pp_2_46_0;
  assign pp_3_46_3 = pp_2_46_1;
  assign pp_3_46_4 = pp_2_46_2;
  assign pp_3_46_5 = pp_2_46_3;
  assign pp_3_46_6 = pp_2_46_4;
  assign pp_3_46_7 = pp_2_46_5;
  assign pp_3_46_8 = pp_2_46_6;
  MG_FA fa_2_47_0(
    .a(pp_2_47_0),
    .b(pp_2_47_1),
    .cin(pp_2_47_2),
    .sum(pp_3_47_0),
    .cout(pp_3_48_0)
  );

  assign pp_3_47_1 = pp_2_47_3;
  assign pp_3_47_2 = pp_2_47_4;
  assign pp_3_48_1 = pp_2_48_0;
  assign pp_3_48_2 = pp_2_48_1;
  assign pp_3_48_3 = pp_2_48_2;
  assign pp_3_48_4 = pp_2_48_3;
  assign pp_3_48_5 = pp_2_48_4;
  MG_FA fa_2_49_0(
    .a(pp_2_49_0),
    .b(pp_2_49_1),
    .cin(pp_2_49_2),
    .sum(pp_3_49_0),
    .cout(pp_3_50_0)
  );

  MG_FA fa_2_49_1(
    .a(pp_2_49_3),
    .b(pp_2_49_4),
    .cin(pp_2_49_5),
    .sum(pp_3_49_1),
    .cout(pp_3_50_1)
  );

  MG_FA fa_2_50_0(
    .a(pp_2_50_0),
    .b(pp_2_50_1),
    .cin(pp_2_50_2),
    .sum(pp_3_50_2),
    .cout(pp_3_51_0)
  );

  MG_FA fa_2_51_0(
    .a(pp_2_51_0),
    .b(pp_2_51_1),
    .cin(pp_2_51_2),
    .sum(pp_3_51_1),
    .cout(pp_3_52_0)
  );

  assign pp_3_51_2 = pp_2_51_3;
  assign pp_3_51_3 = pp_2_51_4;
  MG_FA fa_2_52_0(
    .a(pp_2_52_0),
    .b(pp_2_52_1),
    .cin(pp_2_52_2),
    .sum(pp_3_52_1),
    .cout(pp_3_53_0)
  );

  assign pp_3_52_2 = pp_2_52_3;
  MG_FA fa_2_53_0(
    .a(pp_2_53_0),
    .b(pp_2_53_1),
    .cin(pp_2_53_2),
    .sum(pp_3_53_1),
    .cout(pp_3_54_0)
  );

  assign pp_3_53_2 = pp_2_53_3;
  assign pp_3_53_3 = pp_2_53_4;
  assign pp_3_54_1 = pp_2_54_0;
  assign pp_3_54_2 = pp_2_54_1;
  assign pp_3_54_3 = pp_2_54_2;
  assign pp_3_54_4 = pp_2_54_3;
  MG_FA fa_2_55_0(
    .a(pp_2_55_0),
    .b(pp_2_55_1),
    .cin(pp_2_55_2),
    .sum(pp_3_55_0),
    .cout(pp_3_56_0)
  );

  assign pp_3_55_1 = pp_2_55_3;
  assign pp_3_55_2 = pp_2_55_4;
  MG_FA fa_2_56_0(
    .a(pp_2_56_0),
    .b(pp_2_56_1),
    .cin(pp_2_56_2),
    .sum(pp_3_56_1),
    .cout(pp_3_57_0)
  );

  MG_FA fa_2_56_1(
    .a(pp_2_56_3),
    .b(pp_2_56_4),
    .cin(pp_2_56_5),
    .sum(pp_3_56_2),
    .cout(pp_3_57_1)
  );

  assign pp_3_57_2 = pp_2_57_0;
  assign pp_3_57_3 = pp_2_57_1;
  assign pp_3_58_0 = pp_2_58_0;
  assign pp_3_58_1 = pp_2_58_1;
  assign pp_3_58_2 = pp_2_58_2;
  assign pp_3_59_0 = pp_2_59_0;
  assign pp_3_59_1 = pp_2_59_1;
  assign pp_3_59_2 = pp_2_59_2;
  assign pp_3_59_3 = pp_2_59_3;
  assign pp_3_60_0 = pp_2_60_0;
  MG_FA fa_2_61_0(
    .a(pp_2_61_0),
    .b(pp_2_61_1),
    .cin(pp_2_61_2),
    .sum(pp_3_61_0),
    .cout(pp_3_62_0)
  );

  assign pp_3_62_1 = pp_2_62_0;
  assign pp_3_62_2 = pp_2_62_1;
  MG_FA fa_2_63_0(
    .a(pp_2_63_0),
    .b(pp_2_63_1),
    .cin(pp_2_63_2),
    .sum(pp_3_63_0),
    .cout()
  );

  assign pp_4_0_0 = pp_3_0_0;
  assign pp_4_0_1 = pp_3_0_1;
  assign pp_4_1_0 = pp_3_1_0;
  assign pp_4_2_0 = pp_3_2_0;
  assign pp_4_2_1 = pp_3_2_1;
  assign pp_4_3_0 = pp_3_3_0;
  assign pp_4_3_1 = pp_3_3_1;
  assign pp_4_4_0 = pp_3_4_0;
  assign pp_4_4_1 = pp_3_4_1;
  assign pp_4_4_2 = pp_3_4_2;
  assign pp_4_5_0 = pp_3_5_0;
  assign pp_4_6_0 = pp_3_6_0;
  assign pp_4_6_1 = pp_3_6_1;
  assign pp_4_6_2 = pp_3_6_2;
  assign pp_4_7_0 = pp_3_7_0;
  assign pp_4_8_0 = pp_3_8_0;
  assign pp_4_8_1 = pp_3_8_1;
  assign pp_4_8_2 = pp_3_8_2;
  MG_FA fa_3_9_0(
    .a(pp_3_9_0),
    .b(pp_3_9_1),
    .cin(pp_3_9_2),
    .sum(pp_4_9_0),
    .cout(pp_4_10_0)
  );

  assign pp_4_9_1 = pp_3_9_3;
  assign pp_4_10_1 = pp_3_10_0;
  MG_HA ha_3_11_0(
    .a(pp_3_11_0),
    .b(pp_3_11_1),
    .sum(pp_4_11_0),
    .cout(pp_4_12_0)
  );

  MG_HA ha_3_12_0(
    .a(pp_3_12_0),
    .b(pp_3_12_1),
    .sum(pp_4_12_1),
    .cout(pp_4_13_0)
  );

  MG_FA fa_3_13_0(
    .a(pp_3_13_0),
    .b(pp_3_13_1),
    .cin(pp_3_13_2),
    .sum(pp_4_13_1),
    .cout(pp_4_14_0)
  );

  assign pp_4_13_2 = pp_3_13_3;
  MG_FA fa_3_14_0(
    .a(pp_3_14_0),
    .b(pp_3_14_1),
    .cin(pp_3_14_2),
    .sum(pp_4_14_1),
    .cout(pp_4_15_0)
  );

  MG_FA fa_3_15_0(
    .a(pp_3_15_0),
    .b(pp_3_15_1),
    .cin(pp_3_15_2),
    .sum(pp_4_15_1),
    .cout(pp_4_16_0)
  );

  MG_FA fa_3_16_0(
    .a(pp_3_16_0),
    .b(pp_3_16_1),
    .cin(pp_3_16_2),
    .sum(pp_4_16_1),
    .cout(pp_4_17_0)
  );

  assign pp_4_16_2 = pp_3_16_3;
  MG_FA fa_3_17_0(
    .a(pp_3_17_0),
    .b(pp_3_17_1),
    .cin(pp_3_17_2),
    .sum(pp_4_17_1),
    .cout(pp_4_18_0)
  );

  MG_FA fa_3_18_0(
    .a(pp_3_18_0),
    .b(pp_3_18_1),
    .cin(pp_3_18_2),
    .sum(pp_4_18_1),
    .cout(pp_4_19_0)
  );

  MG_FA fa_3_19_0(
    .a(pp_3_19_0),
    .b(pp_3_19_1),
    .cin(pp_3_19_2),
    .sum(pp_4_19_1),
    .cout(pp_4_20_0)
  );

  assign pp_4_19_2 = pp_3_19_3;
  MG_FA fa_3_20_0(
    .a(pp_3_20_0),
    .b(pp_3_20_1),
    .cin(pp_3_20_2),
    .sum(pp_4_20_1),
    .cout(pp_4_21_0)
  );

  assign pp_4_20_2 = pp_3_20_3;
  MG_FA fa_3_21_0(
    .a(pp_3_21_0),
    .b(pp_3_21_1),
    .cin(pp_3_21_2),
    .sum(pp_4_21_1),
    .cout(pp_4_22_0)
  );

  assign pp_4_21_2 = pp_3_21_3;
  MG_FA fa_3_22_0(
    .a(pp_3_22_0),
    .b(pp_3_22_1),
    .cin(pp_3_22_2),
    .sum(pp_4_22_1),
    .cout(pp_4_23_0)
  );

  MG_FA fa_3_22_1(
    .a(pp_3_22_3),
    .b(pp_3_22_4),
    .cin(pp_3_22_5),
    .sum(pp_4_22_2),
    .cout(pp_4_23_1)
  );

  MG_FA fa_3_23_0(
    .a(pp_3_23_0),
    .b(pp_3_23_1),
    .cin(pp_3_23_2),
    .sum(pp_4_23_2),
    .cout(pp_4_24_0)
  );

  assign pp_4_23_3 = pp_3_23_3;
  MG_FA fa_3_24_0(
    .a(pp_3_24_0),
    .b(pp_3_24_1),
    .cin(pp_3_24_2),
    .sum(pp_4_24_1),
    .cout(pp_4_25_0)
  );

  MG_FA fa_3_24_1(
    .a(pp_3_24_3),
    .b(pp_3_24_4),
    .cin(pp_3_24_5),
    .sum(pp_4_24_2),
    .cout(pp_4_25_1)
  );

  MG_FA fa_3_25_0(
    .a(pp_3_25_0),
    .b(pp_3_25_1),
    .cin(pp_3_25_2),
    .sum(pp_4_25_2),
    .cout(pp_4_26_0)
  );

  MG_FA fa_3_25_1(
    .a(pp_3_25_3),
    .b(pp_3_25_4),
    .cin(pp_3_25_5),
    .sum(pp_4_25_3),
    .cout(pp_4_26_1)
  );

  MG_FA fa_3_26_0(
    .a(pp_3_26_0),
    .b(pp_3_26_1),
    .cin(pp_3_26_2),
    .sum(pp_4_26_2),
    .cout(pp_4_27_0)
  );

  MG_FA fa_3_27_0(
    .a(pp_3_27_0),
    .b(pp_3_27_1),
    .cin(pp_3_27_2),
    .sum(pp_4_27_1),
    .cout(pp_4_28_0)
  );

  MG_FA fa_3_27_1(
    .a(pp_3_27_3),
    .b(pp_3_27_4),
    .cin(pp_3_27_5),
    .sum(pp_4_27_2),
    .cout(pp_4_28_1)
  );

  MG_HA ha_3_28_0(
    .a(pp_3_28_0),
    .b(pp_3_28_1),
    .sum(pp_4_28_2),
    .cout(pp_4_29_0)
  );

  assign pp_4_28_3 = pp_3_28_2;
  assign pp_4_28_4 = pp_3_28_3;
  assign pp_4_28_5 = pp_3_28_4;
  MG_FA fa_3_29_0(
    .a(pp_3_29_0),
    .b(pp_3_29_1),
    .cin(pp_3_29_2),
    .sum(pp_4_29_1),
    .cout(pp_4_30_0)
  );

  MG_HA ha_3_29_1(
    .a(pp_3_29_3),
    .b(pp_3_29_4),
    .sum(pp_4_29_2),
    .cout(pp_4_30_1)
  );

  MG_FA fa_3_30_0(
    .a(pp_3_30_0),
    .b(pp_3_30_1),
    .cin(pp_3_30_2),
    .sum(pp_4_30_2),
    .cout(pp_4_31_0)
  );

  MG_FA fa_3_30_1(
    .a(pp_3_30_3),
    .b(pp_3_30_4),
    .cin(pp_3_30_5),
    .sum(pp_4_30_3),
    .cout(pp_4_31_1)
  );

  MG_FA fa_3_31_0(
    .a(pp_3_31_0),
    .b(pp_3_31_1),
    .cin(pp_3_31_2),
    .sum(pp_4_31_2),
    .cout(pp_4_32_0)
  );

  assign pp_4_31_3 = pp_3_31_3;
  assign pp_4_31_4 = pp_3_31_4;
  assign pp_4_31_5 = pp_3_31_5;
  MG_FA fa_3_32_0(
    .a(pp_3_32_0),
    .b(pp_3_32_1),
    .cin(pp_3_32_2),
    .sum(pp_4_32_1),
    .cout(pp_4_33_0)
  );

  MG_FA fa_3_32_1(
    .a(pp_3_32_3),
    .b(pp_3_32_4),
    .cin(pp_3_32_5),
    .sum(pp_4_32_2),
    .cout(pp_4_33_1)
  );

  MG_FA fa_3_33_0(
    .a(pp_3_33_0),
    .b(pp_3_33_1),
    .cin(pp_3_33_2),
    .sum(pp_4_33_2),
    .cout(pp_4_34_0)
  );

  MG_FA fa_3_33_1(
    .a(pp_3_33_3),
    .b(pp_3_33_4),
    .cin(pp_3_33_5),
    .sum(pp_4_33_3),
    .cout(pp_4_34_1)
  );

  MG_FA fa_3_34_0(
    .a(pp_3_34_0),
    .b(pp_3_34_1),
    .cin(pp_3_34_2),
    .sum(pp_4_34_2),
    .cout(pp_4_35_0)
  );

  MG_FA fa_3_34_1(
    .a(pp_3_34_3),
    .b(pp_3_34_4),
    .cin(pp_3_34_5),
    .sum(pp_4_34_3),
    .cout(pp_4_35_1)
  );

  MG_FA fa_3_35_0(
    .a(pp_3_35_0),
    .b(pp_3_35_1),
    .cin(pp_3_35_2),
    .sum(pp_4_35_2),
    .cout(pp_4_36_0)
  );

  MG_FA fa_3_35_1(
    .a(pp_3_35_3),
    .b(pp_3_35_4),
    .cin(pp_3_35_5),
    .sum(pp_4_35_3),
    .cout(pp_4_36_1)
  );

  MG_FA fa_3_36_0(
    .a(pp_3_36_0),
    .b(pp_3_36_1),
    .cin(pp_3_36_2),
    .sum(pp_4_36_2),
    .cout(pp_4_37_0)
  );

  assign pp_4_36_3 = pp_3_36_3;
  assign pp_4_36_4 = pp_3_36_4;
  MG_FA fa_3_37_0(
    .a(pp_3_37_0),
    .b(pp_3_37_1),
    .cin(pp_3_37_2),
    .sum(pp_4_37_1),
    .cout(pp_4_38_0)
  );

  MG_FA fa_3_37_1(
    .a(pp_3_37_3),
    .b(pp_3_37_4),
    .cin(pp_3_37_5),
    .sum(pp_4_37_2),
    .cout(pp_4_38_1)
  );

  MG_FA fa_3_38_0(
    .a(pp_3_38_0),
    .b(pp_3_38_1),
    .cin(pp_3_38_2),
    .sum(pp_4_38_2),
    .cout(pp_4_39_0)
  );

  MG_FA fa_3_38_1(
    .a(pp_3_38_3),
    .b(pp_3_38_4),
    .cin(pp_3_38_5),
    .sum(pp_4_38_3),
    .cout(pp_4_39_1)
  );

  MG_FA fa_3_39_0(
    .a(pp_3_39_0),
    .b(pp_3_39_1),
    .cin(pp_3_39_2),
    .sum(pp_4_39_2),
    .cout(pp_4_40_0)
  );

  MG_FA fa_3_39_1(
    .a(pp_3_39_3),
    .b(pp_3_39_4),
    .cin(pp_3_39_5),
    .sum(pp_4_39_3),
    .cout(pp_4_40_1)
  );

  MG_HA ha_3_40_0(
    .a(pp_3_40_0),
    .b(pp_3_40_1),
    .sum(pp_4_40_2),
    .cout(pp_4_41_0)
  );

  assign pp_4_40_3 = pp_3_40_2;
  assign pp_4_40_4 = pp_3_40_3;
  assign pp_4_40_5 = pp_3_40_4;
  MG_FA fa_3_41_0(
    .a(pp_3_41_0),
    .b(pp_3_41_1),
    .cin(pp_3_41_2),
    .sum(pp_4_41_1),
    .cout(pp_4_42_0)
  );

  MG_FA fa_3_41_1(
    .a(pp_3_41_3),
    .b(pp_3_41_4),
    .cin(pp_3_41_5),
    .sum(pp_4_41_2),
    .cout(pp_4_42_1)
  );

  MG_FA fa_3_42_0(
    .a(pp_3_42_0),
    .b(pp_3_42_1),
    .cin(pp_3_42_2),
    .sum(pp_4_42_2),
    .cout(pp_4_43_0)
  );

  MG_FA fa_3_43_0(
    .a(pp_3_43_0),
    .b(pp_3_43_1),
    .cin(pp_3_43_2),
    .sum(pp_4_43_1),
    .cout(pp_4_44_0)
  );

  assign pp_4_43_2 = pp_3_43_3;
  assign pp_4_43_3 = pp_3_43_4;
  MG_FA fa_3_44_0(
    .a(pp_3_44_0),
    .b(pp_3_44_1),
    .cin(pp_3_44_2),
    .sum(pp_4_44_1),
    .cout(pp_4_45_0)
  );

  MG_FA fa_3_44_1(
    .a(pp_3_44_3),
    .b(pp_3_44_4),
    .cin(pp_3_44_5),
    .sum(pp_4_44_2),
    .cout(pp_4_45_1)
  );

  assign pp_4_45_2 = pp_3_45_0;
  assign pp_4_45_3 = pp_3_45_1;
  assign pp_4_45_4 = pp_3_45_2;
  assign pp_4_45_5 = pp_3_45_3;
  MG_FA fa_3_46_0(
    .a(pp_3_46_0),
    .b(pp_3_46_1),
    .cin(pp_3_46_2),
    .sum(pp_4_46_0),
    .cout(pp_4_47_0)
  );

  MG_FA fa_3_46_1(
    .a(pp_3_46_3),
    .b(pp_3_46_4),
    .cin(pp_3_46_5),
    .sum(pp_4_46_1),
    .cout(pp_4_47_1)
  );

  MG_FA fa_3_46_2(
    .a(pp_3_46_6),
    .b(pp_3_46_7),
    .cin(pp_3_46_8),
    .sum(pp_4_46_2),
    .cout(pp_4_47_2)
  );

  assign pp_4_47_3 = pp_3_47_0;
  assign pp_4_47_4 = pp_3_47_1;
  assign pp_4_47_5 = pp_3_47_2;
  MG_FA fa_3_48_0(
    .a(pp_3_48_0),
    .b(pp_3_48_1),
    .cin(pp_3_48_2),
    .sum(pp_4_48_0),
    .cout(pp_4_49_0)
  );

  MG_FA fa_3_48_1(
    .a(pp_3_48_3),
    .b(pp_3_48_4),
    .cin(pp_3_48_5),
    .sum(pp_4_48_1),
    .cout(pp_4_49_1)
  );

  assign pp_4_49_2 = pp_3_49_0;
  assign pp_4_49_3 = pp_3_49_1;
  MG_FA fa_3_50_0(
    .a(pp_3_50_0),
    .b(pp_3_50_1),
    .cin(pp_3_50_2),
    .sum(pp_4_50_0),
    .cout(pp_4_51_0)
  );

  MG_FA fa_3_51_0(
    .a(pp_3_51_0),
    .b(pp_3_51_1),
    .cin(pp_3_51_2),
    .sum(pp_4_51_1),
    .cout(pp_4_52_0)
  );

  assign pp_4_51_2 = pp_3_51_3;
  MG_FA fa_3_52_0(
    .a(pp_3_52_0),
    .b(pp_3_52_1),
    .cin(pp_3_52_2),
    .sum(pp_4_52_1),
    .cout(pp_4_53_0)
  );

  MG_FA fa_3_53_0(
    .a(pp_3_53_0),
    .b(pp_3_53_1),
    .cin(pp_3_53_2),
    .sum(pp_4_53_1),
    .cout(pp_4_54_0)
  );

  assign pp_4_53_2 = pp_3_53_3;
  assign pp_4_54_1 = pp_3_54_0;
  assign pp_4_54_2 = pp_3_54_1;
  assign pp_4_54_3 = pp_3_54_2;
  assign pp_4_54_4 = pp_3_54_3;
  assign pp_4_54_5 = pp_3_54_4;
  MG_FA fa_3_55_0(
    .a(pp_3_55_0),
    .b(pp_3_55_1),
    .cin(pp_3_55_2),
    .sum(pp_4_55_0),
    .cout(pp_4_56_0)
  );

  MG_FA fa_3_56_0(
    .a(pp_3_56_0),
    .b(pp_3_56_1),
    .cin(pp_3_56_2),
    .sum(pp_4_56_1),
    .cout(pp_4_57_0)
  );

  MG_FA fa_3_57_0(
    .a(pp_3_57_0),
    .b(pp_3_57_1),
    .cin(pp_3_57_2),
    .sum(pp_4_57_1),
    .cout(pp_4_58_0)
  );

  assign pp_4_57_2 = pp_3_57_3;
  MG_FA fa_3_58_0(
    .a(pp_3_58_0),
    .b(pp_3_58_1),
    .cin(pp_3_58_2),
    .sum(pp_4_58_1),
    .cout(pp_4_59_0)
  );

  MG_FA fa_3_59_0(
    .a(pp_3_59_0),
    .b(pp_3_59_1),
    .cin(pp_3_59_2),
    .sum(pp_4_59_1),
    .cout(pp_4_60_0)
  );

  assign pp_4_59_2 = pp_3_59_3;
  assign pp_4_60_1 = pp_3_60_0;
  assign pp_4_61_0 = pp_3_61_0;
  assign pp_4_62_0 = pp_3_62_0;
  assign pp_4_62_1 = pp_3_62_1;
  assign pp_4_62_2 = pp_3_62_2;
  assign pp_4_63_0 = pp_3_63_0;
  assign pp_5_0_0 = pp_4_0_0;
  assign pp_5_0_1 = pp_4_0_1;
  assign pp_5_1_0 = pp_4_1_0;
  assign pp_5_2_0 = pp_4_2_0;
  assign pp_5_2_1 = pp_4_2_1;
  assign pp_5_3_0 = pp_4_3_0;
  assign pp_5_3_1 = pp_4_3_1;
  MG_HA ha_4_4_0(
    .a(pp_4_4_0),
    .b(pp_4_4_1),
    .sum(pp_5_4_0),
    .cout(pp_5_5_0)
  );

  assign pp_5_4_1 = pp_4_4_2;
  assign pp_5_5_1 = pp_4_5_0;
  MG_HA ha_4_6_0(
    .a(pp_4_6_0),
    .b(pp_4_6_1),
    .sum(pp_5_6_0),
    .cout(pp_5_7_0)
  );

  assign pp_5_6_1 = pp_4_6_2;
  assign pp_5_7_1 = pp_4_7_0;
  assign pp_5_8_0 = pp_4_8_0;
  assign pp_5_8_1 = pp_4_8_1;
  assign pp_5_8_2 = pp_4_8_2;
  MG_HA ha_4_9_0(
    .a(pp_4_9_0),
    .b(pp_4_9_1),
    .sum(pp_5_9_0),
    .cout(pp_5_10_0)
  );

  MG_HA ha_4_10_0(
    .a(pp_4_10_0),
    .b(pp_4_10_1),
    .sum(pp_5_10_1),
    .cout(pp_5_11_0)
  );

  assign pp_5_11_1 = pp_4_11_0;
  assign pp_5_12_0 = pp_4_12_0;
  assign pp_5_12_1 = pp_4_12_1;
  assign pp_5_13_0 = pp_4_13_0;
  assign pp_5_13_1 = pp_4_13_1;
  assign pp_5_13_2 = pp_4_13_2;
  MG_HA ha_4_14_0(
    .a(pp_4_14_0),
    .b(pp_4_14_1),
    .sum(pp_5_14_0),
    .cout(pp_5_15_0)
  );

  assign pp_5_15_1 = pp_4_15_0;
  assign pp_5_15_2 = pp_4_15_1;
  MG_FA fa_4_16_0(
    .a(pp_4_16_0),
    .b(pp_4_16_1),
    .cin(pp_4_16_2),
    .sum(pp_5_16_0),
    .cout(pp_5_17_0)
  );

  assign pp_5_17_1 = pp_4_17_0;
  assign pp_5_17_2 = pp_4_17_1;
  MG_HA ha_4_18_0(
    .a(pp_4_18_0),
    .b(pp_4_18_1),
    .sum(pp_5_18_0),
    .cout(pp_5_19_0)
  );

  assign pp_5_19_1 = pp_4_19_0;
  assign pp_5_19_2 = pp_4_19_1;
  assign pp_5_19_3 = pp_4_19_2;
  MG_FA fa_4_20_0(
    .a(pp_4_20_0),
    .b(pp_4_20_1),
    .cin(pp_4_20_2),
    .sum(pp_5_20_0),
    .cout(pp_5_21_0)
  );

  assign pp_5_21_1 = pp_4_21_0;
  assign pp_5_21_2 = pp_4_21_1;
  assign pp_5_21_3 = pp_4_21_2;
  MG_FA fa_4_22_0(
    .a(pp_4_22_0),
    .b(pp_4_22_1),
    .cin(pp_4_22_2),
    .sum(pp_5_22_0),
    .cout(pp_5_23_0)
  );

  MG_HA ha_4_23_0(
    .a(pp_4_23_0),
    .b(pp_4_23_1),
    .sum(pp_5_23_1),
    .cout(pp_5_24_0)
  );

  assign pp_5_23_2 = pp_4_23_2;
  assign pp_5_23_3 = pp_4_23_3;
  MG_HA ha_4_24_0(
    .a(pp_4_24_0),
    .b(pp_4_24_1),
    .sum(pp_5_24_1),
    .cout(pp_5_25_0)
  );

  assign pp_5_24_2 = pp_4_24_2;
  MG_FA fa_4_25_0(
    .a(pp_4_25_0),
    .b(pp_4_25_1),
    .cin(pp_4_25_2),
    .sum(pp_5_25_1),
    .cout(pp_5_26_0)
  );

  assign pp_5_25_2 = pp_4_25_3;
  MG_FA fa_4_26_0(
    .a(pp_4_26_0),
    .b(pp_4_26_1),
    .cin(pp_4_26_2),
    .sum(pp_5_26_1),
    .cout(pp_5_27_0)
  );

  MG_FA fa_4_27_0(
    .a(pp_4_27_0),
    .b(pp_4_27_1),
    .cin(pp_4_27_2),
    .sum(pp_5_27_1),
    .cout(pp_5_28_0)
  );

  MG_FA fa_4_28_0(
    .a(pp_4_28_0),
    .b(pp_4_28_1),
    .cin(pp_4_28_2),
    .sum(pp_5_28_1),
    .cout(pp_5_29_0)
  );

  MG_FA fa_4_28_1(
    .a(pp_4_28_3),
    .b(pp_4_28_4),
    .cin(pp_4_28_5),
    .sum(pp_5_28_2),
    .cout(pp_5_29_1)
  );

  MG_FA fa_4_29_0(
    .a(pp_4_29_0),
    .b(pp_4_29_1),
    .cin(pp_4_29_2),
    .sum(pp_5_29_2),
    .cout(pp_5_30_0)
  );

  MG_FA fa_4_30_0(
    .a(pp_4_30_0),
    .b(pp_4_30_1),
    .cin(pp_4_30_2),
    .sum(pp_5_30_1),
    .cout(pp_5_31_0)
  );

  assign pp_5_30_2 = pp_4_30_3;
  MG_FA fa_4_31_0(
    .a(pp_4_31_0),
    .b(pp_4_31_1),
    .cin(pp_4_31_2),
    .sum(pp_5_31_1),
    .cout(pp_5_32_0)
  );

  MG_FA fa_4_31_1(
    .a(pp_4_31_3),
    .b(pp_4_31_4),
    .cin(pp_4_31_5),
    .sum(pp_5_31_2),
    .cout(pp_5_32_1)
  );

  MG_FA fa_4_32_0(
    .a(pp_4_32_0),
    .b(pp_4_32_1),
    .cin(pp_4_32_2),
    .sum(pp_5_32_2),
    .cout(pp_5_33_0)
  );

  MG_FA fa_4_33_0(
    .a(pp_4_33_0),
    .b(pp_4_33_1),
    .cin(pp_4_33_2),
    .sum(pp_5_33_1),
    .cout(pp_5_34_0)
  );

  assign pp_5_33_2 = pp_4_33_3;
  MG_FA fa_4_34_0(
    .a(pp_4_34_0),
    .b(pp_4_34_1),
    .cin(pp_4_34_2),
    .sum(pp_5_34_1),
    .cout(pp_5_35_0)
  );

  assign pp_5_34_2 = pp_4_34_3;
  MG_FA fa_4_35_0(
    .a(pp_4_35_0),
    .b(pp_4_35_1),
    .cin(pp_4_35_2),
    .sum(pp_5_35_1),
    .cout(pp_5_36_0)
  );

  assign pp_5_35_2 = pp_4_35_3;
  MG_FA fa_4_36_0(
    .a(pp_4_36_0),
    .b(pp_4_36_1),
    .cin(pp_4_36_2),
    .sum(pp_5_36_1),
    .cout(pp_5_37_0)
  );

  MG_HA ha_4_36_1(
    .a(pp_4_36_3),
    .b(pp_4_36_4),
    .sum(pp_5_36_2),
    .cout(pp_5_37_1)
  );

  MG_FA fa_4_37_0(
    .a(pp_4_37_0),
    .b(pp_4_37_1),
    .cin(pp_4_37_2),
    .sum(pp_5_37_2),
    .cout(pp_5_38_0)
  );

  MG_FA fa_4_38_0(
    .a(pp_4_38_0),
    .b(pp_4_38_1),
    .cin(pp_4_38_2),
    .sum(pp_5_38_1),
    .cout(pp_5_39_0)
  );

  assign pp_5_38_2 = pp_4_38_3;
  MG_FA fa_4_39_0(
    .a(pp_4_39_0),
    .b(pp_4_39_1),
    .cin(pp_4_39_2),
    .sum(pp_5_39_1),
    .cout(pp_5_40_0)
  );

  assign pp_5_39_2 = pp_4_39_3;
  MG_FA fa_4_40_0(
    .a(pp_4_40_0),
    .b(pp_4_40_1),
    .cin(pp_4_40_2),
    .sum(pp_5_40_1),
    .cout(pp_5_41_0)
  );

  MG_FA fa_4_40_1(
    .a(pp_4_40_3),
    .b(pp_4_40_4),
    .cin(pp_4_40_5),
    .sum(pp_5_40_2),
    .cout(pp_5_41_1)
  );

  MG_FA fa_4_41_0(
    .a(pp_4_41_0),
    .b(pp_4_41_1),
    .cin(pp_4_41_2),
    .sum(pp_5_41_2),
    .cout(pp_5_42_0)
  );

  MG_HA ha_4_42_0(
    .a(pp_4_42_0),
    .b(pp_4_42_1),
    .sum(pp_5_42_1),
    .cout(pp_5_43_0)
  );

  assign pp_5_42_2 = pp_4_42_2;
  MG_FA fa_4_43_0(
    .a(pp_4_43_0),
    .b(pp_4_43_1),
    .cin(pp_4_43_2),
    .sum(pp_5_43_1),
    .cout(pp_5_44_0)
  );

  assign pp_5_43_2 = pp_4_43_3;
  MG_FA fa_4_44_0(
    .a(pp_4_44_0),
    .b(pp_4_44_1),
    .cin(pp_4_44_2),
    .sum(pp_5_44_1),
    .cout(pp_5_45_0)
  );

  MG_FA fa_4_45_0(
    .a(pp_4_45_0),
    .b(pp_4_45_1),
    .cin(pp_4_45_2),
    .sum(pp_5_45_1),
    .cout(pp_5_46_0)
  );

  MG_FA fa_4_45_1(
    .a(pp_4_45_3),
    .b(pp_4_45_4),
    .cin(pp_4_45_5),
    .sum(pp_5_45_2),
    .cout(pp_5_46_1)
  );

  MG_FA fa_4_46_0(
    .a(pp_4_46_0),
    .b(pp_4_46_1),
    .cin(pp_4_46_2),
    .sum(pp_5_46_2),
    .cout(pp_5_47_0)
  );

  MG_FA fa_4_47_0(
    .a(pp_4_47_0),
    .b(pp_4_47_1),
    .cin(pp_4_47_2),
    .sum(pp_5_47_1),
    .cout(pp_5_48_0)
  );

  MG_FA fa_4_47_1(
    .a(pp_4_47_3),
    .b(pp_4_47_4),
    .cin(pp_4_47_5),
    .sum(pp_5_47_2),
    .cout(pp_5_48_1)
  );

  MG_HA ha_4_48_0(
    .a(pp_4_48_0),
    .b(pp_4_48_1),
    .sum(pp_5_48_2),
    .cout(pp_5_49_0)
  );

  MG_FA fa_4_49_0(
    .a(pp_4_49_0),
    .b(pp_4_49_1),
    .cin(pp_4_49_2),
    .sum(pp_5_49_1),
    .cout(pp_5_50_0)
  );

  assign pp_5_49_2 = pp_4_49_3;
  assign pp_5_50_1 = pp_4_50_0;
  assign pp_5_51_0 = pp_4_51_0;
  assign pp_5_51_1 = pp_4_51_1;
  assign pp_5_51_2 = pp_4_51_2;
  MG_HA ha_4_52_0(
    .a(pp_4_52_0),
    .b(pp_4_52_1),
    .sum(pp_5_52_0),
    .cout(pp_5_53_0)
  );

  assign pp_5_53_1 = pp_4_53_0;
  assign pp_5_53_2 = pp_4_53_1;
  assign pp_5_53_3 = pp_4_53_2;
  MG_FA fa_4_54_0(
    .a(pp_4_54_0),
    .b(pp_4_54_1),
    .cin(pp_4_54_2),
    .sum(pp_5_54_0),
    .cout(pp_5_55_0)
  );

  MG_FA fa_4_54_1(
    .a(pp_4_54_3),
    .b(pp_4_54_4),
    .cin(pp_4_54_5),
    .sum(pp_5_54_1),
    .cout(pp_5_55_1)
  );

  assign pp_5_55_2 = pp_4_55_0;
  assign pp_5_56_0 = pp_4_56_0;
  assign pp_5_56_1 = pp_4_56_1;
  assign pp_5_57_0 = pp_4_57_0;
  assign pp_5_57_1 = pp_4_57_1;
  assign pp_5_57_2 = pp_4_57_2;
  assign pp_5_58_0 = pp_4_58_0;
  assign pp_5_58_1 = pp_4_58_1;
  MG_FA fa_4_59_0(
    .a(pp_4_59_0),
    .b(pp_4_59_1),
    .cin(pp_4_59_2),
    .sum(pp_5_59_0),
    .cout(pp_5_60_0)
  );

  assign pp_5_60_1 = pp_4_60_0;
  assign pp_5_60_2 = pp_4_60_1;
  assign pp_5_61_0 = pp_4_61_0;
  assign pp_5_62_0 = pp_4_62_0;
  assign pp_5_62_1 = pp_4_62_1;
  assign pp_5_62_2 = pp_4_62_2;
  assign pp_5_63_0 = pp_4_63_0;
  assign pp_6_0_0 = pp_5_0_0;
  assign pp_6_0_1 = pp_5_0_1;
  assign pp_6_1_0 = pp_5_1_0;
  assign pp_6_2_0 = pp_5_2_0;
  assign pp_6_2_1 = pp_5_2_1;
  assign pp_6_3_0 = pp_5_3_0;
  assign pp_6_3_1 = pp_5_3_1;
  assign pp_6_4_0 = pp_5_4_0;
  assign pp_6_4_1 = pp_5_4_1;
  assign pp_6_5_0 = pp_5_5_0;
  assign pp_6_5_1 = pp_5_5_1;
  assign pp_6_6_0 = pp_5_6_0;
  assign pp_6_6_1 = pp_5_6_1;
  assign pp_6_7_0 = pp_5_7_0;
  assign pp_6_7_1 = pp_5_7_1;
  MG_HA ha_5_8_0(
    .a(pp_5_8_0),
    .b(pp_5_8_1),
    .sum(pp_6_8_0),
    .cout(pp_6_9_0)
  );

  assign pp_6_8_1 = pp_5_8_2;
  assign pp_6_9_1 = pp_5_9_0;
  assign pp_6_10_0 = pp_5_10_0;
  assign pp_6_10_1 = pp_5_10_1;
  assign pp_6_11_0 = pp_5_11_0;
  assign pp_6_11_1 = pp_5_11_1;
  assign pp_6_12_0 = pp_5_12_0;
  assign pp_6_12_1 = pp_5_12_1;
  MG_HA ha_5_13_0(
    .a(pp_5_13_0),
    .b(pp_5_13_1),
    .sum(pp_6_13_0),
    .cout(pp_6_14_0)
  );

  assign pp_6_13_1 = pp_5_13_2;
  assign pp_6_14_1 = pp_5_14_0;
  MG_HA ha_5_15_0(
    .a(pp_5_15_0),
    .b(pp_5_15_1),
    .sum(pp_6_15_0),
    .cout(pp_6_16_0)
  );

  assign pp_6_15_1 = pp_5_15_2;
  assign pp_6_16_1 = pp_5_16_0;
  MG_HA ha_5_17_0(
    .a(pp_5_17_0),
    .b(pp_5_17_1),
    .sum(pp_6_17_0),
    .cout(pp_6_18_0)
  );

  assign pp_6_17_1 = pp_5_17_2;
  assign pp_6_18_1 = pp_5_18_0;
  MG_FA fa_5_19_0(
    .a(pp_5_19_0),
    .b(pp_5_19_1),
    .cin(pp_5_19_2),
    .sum(pp_6_19_0),
    .cout(pp_6_20_0)
  );

  assign pp_6_19_1 = pp_5_19_3;
  assign pp_6_20_1 = pp_5_20_0;
  MG_FA fa_5_21_0(
    .a(pp_5_21_0),
    .b(pp_5_21_1),
    .cin(pp_5_21_2),
    .sum(pp_6_21_0),
    .cout(pp_6_22_0)
  );

  assign pp_6_21_1 = pp_5_21_3;
  assign pp_6_22_1 = pp_5_22_0;
  MG_FA fa_5_23_0(
    .a(pp_5_23_0),
    .b(pp_5_23_1),
    .cin(pp_5_23_2),
    .sum(pp_6_23_0),
    .cout(pp_6_24_0)
  );

  assign pp_6_23_1 = pp_5_23_3;
  MG_FA fa_5_24_0(
    .a(pp_5_24_0),
    .b(pp_5_24_1),
    .cin(pp_5_24_2),
    .sum(pp_6_24_1),
    .cout(pp_6_25_0)
  );

  MG_FA fa_5_25_0(
    .a(pp_5_25_0),
    .b(pp_5_25_1),
    .cin(pp_5_25_2),
    .sum(pp_6_25_1),
    .cout(pp_6_26_0)
  );

  MG_HA ha_5_26_0(
    .a(pp_5_26_0),
    .b(pp_5_26_1),
    .sum(pp_6_26_1),
    .cout(pp_6_27_0)
  );

  MG_HA ha_5_27_0(
    .a(pp_5_27_0),
    .b(pp_5_27_1),
    .sum(pp_6_27_1),
    .cout(pp_6_28_0)
  );

  MG_FA fa_5_28_0(
    .a(pp_5_28_0),
    .b(pp_5_28_1),
    .cin(pp_5_28_2),
    .sum(pp_6_28_1),
    .cout(pp_6_29_0)
  );

  MG_FA fa_5_29_0(
    .a(pp_5_29_0),
    .b(pp_5_29_1),
    .cin(pp_5_29_2),
    .sum(pp_6_29_1),
    .cout(pp_6_30_0)
  );

  MG_FA fa_5_30_0(
    .a(pp_5_30_0),
    .b(pp_5_30_1),
    .cin(pp_5_30_2),
    .sum(pp_6_30_1),
    .cout(pp_6_31_0)
  );

  MG_FA fa_5_31_0(
    .a(pp_5_31_0),
    .b(pp_5_31_1),
    .cin(pp_5_31_2),
    .sum(pp_6_31_1),
    .cout(pp_6_32_0)
  );

  MG_FA fa_5_32_0(
    .a(pp_5_32_0),
    .b(pp_5_32_1),
    .cin(pp_5_32_2),
    .sum(pp_6_32_1),
    .cout(pp_6_33_0)
  );

  MG_FA fa_5_33_0(
    .a(pp_5_33_0),
    .b(pp_5_33_1),
    .cin(pp_5_33_2),
    .sum(pp_6_33_1),
    .cout(pp_6_34_0)
  );

  MG_FA fa_5_34_0(
    .a(pp_5_34_0),
    .b(pp_5_34_1),
    .cin(pp_5_34_2),
    .sum(pp_6_34_1),
    .cout(pp_6_35_0)
  );

  MG_FA fa_5_35_0(
    .a(pp_5_35_0),
    .b(pp_5_35_1),
    .cin(pp_5_35_2),
    .sum(pp_6_35_1),
    .cout(pp_6_36_0)
  );

  MG_FA fa_5_36_0(
    .a(pp_5_36_0),
    .b(pp_5_36_1),
    .cin(pp_5_36_2),
    .sum(pp_6_36_1),
    .cout(pp_6_37_0)
  );

  MG_FA fa_5_37_0(
    .a(pp_5_37_0),
    .b(pp_5_37_1),
    .cin(pp_5_37_2),
    .sum(pp_6_37_1),
    .cout(pp_6_38_0)
  );

  MG_FA fa_5_38_0(
    .a(pp_5_38_0),
    .b(pp_5_38_1),
    .cin(pp_5_38_2),
    .sum(pp_6_38_1),
    .cout(pp_6_39_0)
  );

  MG_FA fa_5_39_0(
    .a(pp_5_39_0),
    .b(pp_5_39_1),
    .cin(pp_5_39_2),
    .sum(pp_6_39_1),
    .cout(pp_6_40_0)
  );

  MG_FA fa_5_40_0(
    .a(pp_5_40_0),
    .b(pp_5_40_1),
    .cin(pp_5_40_2),
    .sum(pp_6_40_1),
    .cout(pp_6_41_0)
  );

  MG_FA fa_5_41_0(
    .a(pp_5_41_0),
    .b(pp_5_41_1),
    .cin(pp_5_41_2),
    .sum(pp_6_41_1),
    .cout(pp_6_42_0)
  );

  MG_FA fa_5_42_0(
    .a(pp_5_42_0),
    .b(pp_5_42_1),
    .cin(pp_5_42_2),
    .sum(pp_6_42_1),
    .cout(pp_6_43_0)
  );

  MG_FA fa_5_43_0(
    .a(pp_5_43_0),
    .b(pp_5_43_2),
    .cin(pp_5_43_1),
    .sum(pp_6_43_1),
    .cout(pp_6_44_0)
  );

  MG_HA ha_5_44_0(
    .a(pp_5_44_0),
    .b(pp_5_44_1),
    .sum(pp_6_44_1),
    .cout(pp_6_45_0)
  );

  MG_FA fa_5_45_0(
    .a(pp_5_45_0),
    .b(pp_5_45_1),
    .cin(pp_5_45_2),
    .sum(pp_6_45_1),
    .cout(pp_6_46_0)
  );

  MG_FA fa_5_46_0(
    .a(pp_5_46_0),
    .b(pp_5_46_1),
    .cin(pp_5_46_2),
    .sum(pp_6_46_1),
    .cout(pp_6_47_0)
  );

  MG_FA fa_5_47_0(
    .a(pp_5_47_0),
    .b(pp_5_47_1),
    .cin(pp_5_47_2),
    .sum(pp_6_47_1),
    .cout(pp_6_48_0)
  );

  MG_FA fa_5_48_0(
    .a(pp_5_48_0),
    .b(pp_5_48_1),
    .cin(pp_5_48_2),
    .sum(pp_6_48_1),
    .cout(pp_6_49_0)
  );

  MG_FA fa_5_49_0(
    .a(pp_5_49_0),
    .b(pp_5_49_1),
    .cin(pp_5_49_2),
    .sum(pp_6_49_1),
    .cout(pp_6_50_0)
  );

  MG_HA ha_5_50_0(
    .a(pp_5_50_0),
    .b(pp_5_50_1),
    .sum(pp_6_50_1),
    .cout(pp_6_51_0)
  );

  MG_FA fa_5_51_0(
    .a(pp_5_51_0),
    .b(pp_5_51_1),
    .cin(pp_5_51_2),
    .sum(pp_6_51_1),
    .cout(pp_6_52_0)
  );

  assign pp_6_52_1 = pp_5_52_0;
  MG_FA fa_5_53_0(
    .a(pp_5_53_0),
    .b(pp_5_53_1),
    .cin(pp_5_53_2),
    .sum(pp_6_53_0),
    .cout(pp_6_54_0)
  );

  assign pp_6_53_1 = pp_5_53_3;
  MG_HA ha_5_54_0(
    .a(pp_5_54_0),
    .b(pp_5_54_1),
    .sum(pp_6_54_1),
    .cout(pp_6_55_0)
  );

  MG_FA fa_5_55_0(
    .a(pp_5_55_0),
    .b(pp_5_55_1),
    .cin(pp_5_55_2),
    .sum(pp_6_55_1),
    .cout(pp_6_56_0)
  );

  MG_HA ha_5_56_0(
    .a(pp_5_56_0),
    .b(pp_5_56_1),
    .sum(pp_6_56_1),
    .cout(pp_6_57_0)
  );

  MG_FA fa_5_57_0(
    .a(pp_5_57_0),
    .b(pp_5_57_1),
    .cin(pp_5_57_2),
    .sum(pp_6_57_1),
    .cout(pp_6_58_0)
  );

  MG_HA ha_5_58_0(
    .a(pp_5_58_0),
    .b(pp_5_58_1),
    .sum(pp_6_58_1),
    .cout(pp_6_59_0)
  );

  assign pp_6_59_1 = pp_5_59_0;
  MG_HA ha_5_60_0(
    .a(pp_5_60_0),
    .b(pp_5_60_1),
    .sum(pp_6_60_0),
    .cout(pp_6_61_0)
  );

  assign pp_6_60_1 = pp_5_60_2;
  assign pp_6_61_1 = pp_5_61_0;
  MG_HA ha_5_62_0(
    .a(pp_5_62_0),
    .b(pp_5_62_1),
    .sum(pp_6_62_0),
    .cout(pp_6_63_0)
  );

  assign pp_6_62_1 = pp_5_62_2;
  assign pp_6_63_1 = pp_5_63_0;
  wire [63:0] cta;
  wire [63:0] ctb;
  wire [63:0] cts;
  wire ctc;

  MG_CPA cpa(
 .a(cta), .b(ctb), .sum(cts), .cout(ctc)
  );

  assign cta[0] = pp_6_0_0;
  assign ctb[0] = pp_6_0_1;
  assign cta[1] = pp_6_1_0;
  assign ctb[1] = 1'b0;
  assign cta[2] = pp_6_2_0;
  assign ctb[2] = pp_6_2_1;
  assign cta[3] = pp_6_3_0;
  assign ctb[3] = pp_6_3_1;
  assign cta[4] = pp_6_4_0;
  assign ctb[4] = pp_6_4_1;
  assign cta[5] = pp_6_5_0;
  assign ctb[5] = pp_6_5_1;
  assign cta[6] = pp_6_6_0;
  assign ctb[6] = pp_6_6_1;
  assign cta[7] = pp_6_7_0;
  assign ctb[7] = pp_6_7_1;
  assign cta[8] = pp_6_8_0;
  assign ctb[8] = pp_6_8_1;
  assign cta[9] = pp_6_9_0;
  assign ctb[9] = pp_6_9_1;
  assign cta[10] = pp_6_10_0;
  assign ctb[10] = pp_6_10_1;
  assign cta[11] = pp_6_11_0;
  assign ctb[11] = pp_6_11_1;
  assign cta[12] = pp_6_12_0;
  assign ctb[12] = pp_6_12_1;
  assign cta[13] = pp_6_13_0;
  assign ctb[13] = pp_6_13_1;
  assign cta[14] = pp_6_14_0;
  assign ctb[14] = pp_6_14_1;
  assign cta[15] = pp_6_15_0;
  assign ctb[15] = pp_6_15_1;
  assign cta[16] = pp_6_16_0;
  assign ctb[16] = pp_6_16_1;
  assign cta[17] = pp_6_17_0;
  assign ctb[17] = pp_6_17_1;
  assign cta[18] = pp_6_18_0;
  assign ctb[18] = pp_6_18_1;
  assign cta[19] = pp_6_19_0;
  assign ctb[19] = pp_6_19_1;
  assign cta[20] = pp_6_20_0;
  assign ctb[20] = pp_6_20_1;
  assign cta[21] = pp_6_21_0;
  assign ctb[21] = pp_6_21_1;
  assign cta[22] = pp_6_22_0;
  assign ctb[22] = pp_6_22_1;
  assign cta[23] = pp_6_23_0;
  assign ctb[23] = pp_6_23_1;
  assign cta[24] = pp_6_24_0;
  assign ctb[24] = pp_6_24_1;
  assign cta[25] = pp_6_25_0;
  assign ctb[25] = pp_6_25_1;
  assign cta[26] = pp_6_26_0;
  assign ctb[26] = pp_6_26_1;
  assign cta[27] = pp_6_27_0;
  assign ctb[27] = pp_6_27_1;
  assign cta[28] = pp_6_28_0;
  assign ctb[28] = pp_6_28_1;
  assign cta[29] = pp_6_29_0;
  assign ctb[29] = pp_6_29_1;
  assign cta[30] = pp_6_30_0;
  assign ctb[30] = pp_6_30_1;
  assign cta[31] = pp_6_31_0;
  assign ctb[31] = pp_6_31_1;
  assign cta[32] = pp_6_32_0;
  assign ctb[32] = pp_6_32_1;
  assign cta[33] = pp_6_33_0;
  assign ctb[33] = pp_6_33_1;
  assign cta[34] = pp_6_34_0;
  assign ctb[34] = pp_6_34_1;
  assign cta[35] = pp_6_35_0;
  assign ctb[35] = pp_6_35_1;
  assign cta[36] = pp_6_36_0;
  assign ctb[36] = pp_6_36_1;
  assign cta[37] = pp_6_37_0;
  assign ctb[37] = pp_6_37_1;
  assign cta[38] = pp_6_38_0;
  assign ctb[38] = pp_6_38_1;
  assign cta[39] = pp_6_39_0;
  assign ctb[39] = pp_6_39_1;
  assign cta[40] = pp_6_40_0;
  assign ctb[40] = pp_6_40_1;
  assign cta[41] = pp_6_41_0;
  assign ctb[41] = pp_6_41_1;
  assign cta[42] = pp_6_42_0;
  assign ctb[42] = pp_6_42_1;
  assign cta[43] = pp_6_43_0;
  assign ctb[43] = pp_6_43_1;
  assign cta[44] = pp_6_44_0;
  assign ctb[44] = pp_6_44_1;
  assign cta[45] = pp_6_45_0;
  assign ctb[45] = pp_6_45_1;
  assign cta[46] = pp_6_46_0;
  assign ctb[46] = pp_6_46_1;
  assign cta[47] = pp_6_47_0;
  assign ctb[47] = pp_6_47_1;
  assign cta[48] = pp_6_48_0;
  assign ctb[48] = pp_6_48_1;
  assign cta[49] = pp_6_49_0;
  assign ctb[49] = pp_6_49_1;
  assign cta[50] = pp_6_50_0;
  assign ctb[50] = pp_6_50_1;
  assign cta[51] = pp_6_51_0;
  assign ctb[51] = pp_6_51_1;
  assign cta[52] = pp_6_52_0;
  assign ctb[52] = pp_6_52_1;
  assign cta[53] = pp_6_53_0;
  assign ctb[53] = pp_6_53_1;
  assign cta[54] = pp_6_54_0;
  assign ctb[54] = pp_6_54_1;
  assign cta[55] = pp_6_55_0;
  assign ctb[55] = pp_6_55_1;
  assign cta[56] = pp_6_56_0;
  assign ctb[56] = pp_6_56_1;
  assign cta[57] = pp_6_57_0;
  assign ctb[57] = pp_6_57_1;
  assign cta[58] = pp_6_58_0;
  assign ctb[58] = pp_6_58_1;
  assign cta[59] = pp_6_59_0;
  assign ctb[59] = pp_6_59_1;
  assign cta[60] = pp_6_60_0;
  assign ctb[60] = pp_6_60_1;
  assign cta[61] = pp_6_61_0;
  assign ctb[61] = pp_6_61_1;
  assign cta[62] = pp_6_62_0;
  assign ctb[62] = pp_6_62_1;
  assign cta[63] = pp_6_63_0;
  assign ctb[63] = pp_6_63_1;
  assign product[63:0] = cts;
endmodule
