module gemm_mac_int8 #(
    parameter integer LANES = 8,
    parameter integer ACC_WIDTH = 32
) (
    input  wire [LANES*8-1:0] a_vec,
    input  wire [LANES*8-1:0] b_vec,
    output reg  signed [ACC_WIDTH-1:0] acc_out
);
  integer i;
  reg signed [ACC_WIDTH-1:0] sum;
  reg signed [7:0] a_i;
  reg signed [7:0] b_i;

  always @(*) begin
    sum = 0;
    for (i = 0; i < LANES; i = i + 1) begin
      a_i = a_vec[(i*8) +: 8];
      b_i = b_vec[(i*8) +: 8];
      sum = sum + (a_i * b_i);
    end
    acc_out = sum;
  end
endmodule


module gemm_mac_int16 #(
    parameter integer LANES = 4,
    parameter integer ACC_WIDTH = 32
) (
    input  wire [LANES*16-1:0] a_vec,
    input  wire [LANES*16-1:0] b_vec,
    output reg  signed [ACC_WIDTH-1:0] acc_out
);
  integer i;
  reg signed [ACC_WIDTH-1:0] sum;
  reg signed [15:0] a_i;
  reg signed [15:0] b_i;

  always @(*) begin
    sum = 0;
    for (i = 0; i < LANES; i = i + 1) begin
      a_i = a_vec[(i*16) +: 16];
      b_i = b_vec[(i*16) +: 16];
      sum = sum + (a_i * b_i);
    end
    acc_out = sum;
  end
endmodule


module gemm_mac_fp16 #(
    parameter integer LANES = 4,
    parameter integer ACC_WIDTH = 32
) (
    input  wire [LANES*16-1:0] a_vec,
    input  wire [LANES*16-1:0] b_vec,
    output reg  signed [ACC_WIDTH-1:0] acc_out
);
  integer i;
  reg signed [ACC_WIDTH-1:0] sum;
  reg signed [15:0] a_i;
  reg signed [15:0] b_i;

  // Phase-3 placeholder: treat fp16 lanes as raw signed-16 values.
  // Swap this block with true IEEE-754 half MAC when fp16 datapath is integrated.
  always @(*) begin
    sum = 0;
    for (i = 0; i < LANES; i = i + 1) begin
      a_i = a_vec[(i*16) +: 16];
      b_i = b_vec[(i*16) +: 16];
      sum = sum + (a_i * b_i);
    end
    acc_out = sum;
  end
endmodule


// Auto-generated by npu/rtlgen/gen.py (v0.1)
module npu_fp16_builtin_l1 (
    input  wire                  clk,
    input  wire                  rst_n,
    input  wire [11:0] mmio_addr,
    input  wire                  mmio_we,
    input  wire [31:0] mmio_wdata,
    output reg  [31:0] mmio_rdata,
    output reg                   irq,
    output reg                   dma_req_valid,
    output reg  [63:0] dma_req_src,
    output reg  [63:0] dma_req_dst,
    output reg  [31:0]           dma_req_bytes,
    input  wire                  dma_req_ready,
    input  wire                  dma_resp_done
,
    output reg  [63:0] cq_mem_addr,
    input  wire [255:0]          cq_mem_rdata
,
    output reg                   m_axi_awvalid,
    input  wire                  m_axi_awready,
    output reg  [63:0] m_axi_awaddr,
    output reg  [7:0]            m_axi_awlen,
    output reg  [2:0]            m_axi_awsize,
    output reg                   m_axi_wvalid,
    input  wire                  m_axi_wready,
    output reg  [255:0] m_axi_wdata,
    output reg  [31:0] m_axi_wstrb,
    output reg                   m_axi_wlast,
    input  wire                  m_axi_bvalid,
    output reg                   m_axi_bready,
    output reg                   m_axi_arvalid,
    input  wire                  m_axi_arready,
    output reg  [63:0] m_axi_araddr,
    output reg  [7:0]            m_axi_arlen,
    output reg  [2:0]            m_axi_arsize,
    input  wire                  m_axi_rvalid,
    output reg                   m_axi_rready,
    input  wire [255:0] m_axi_rdata,
    input  wire                  m_axi_rlast

);

  // Minimal stub: MMIO register block with queue bookkeeping.
  reg [31:0] version;
  reg [31:0] capabilities;
  reg [31:0] status;
  reg [31:0] control;
  reg [31:0] irq_status;
  reg [31:0] irq_enable;
  reg [31:0] cq_base_lo;
  reg [31:0] cq_base_hi;
  reg [31:0] cq_size;
  reg [31:0] cq_head;
  reg [31:0] cq_tail;
  reg [31:0] cq_count;
  reg [255:0] cq_word0;
  reg [7:0]  cq_word0_size;
  reg        cq_pending_ext;
  reg [7:0] last_opcode;
  reg [31:0] last_tag;
  reg [63:0] last_src;
  reg [63:0] last_dst;
  reg [31:0] last_size;
  reg [63:0] last_op_uid;
  reg [63:0] dma_src;
  reg [63:0] dma_dst;
  reg [31:0] dma_size;
  reg        cq_stage_valid;
  reg        dma_pending;
  reg [2:0]  dma_state;
  reg        gemm_pending;
  reg [1:0]  gemm_slot_valid;
  reg [1:0]  gemm_slot_done;
  reg [31:0] gemm_slot_cycles0;
  reg [31:0] gemm_slot_cycles1;
  reg [63:0] gemm_slot_uid0;
  reg [63:0] gemm_slot_uid1;
  reg [63:0] gemm_slot_src0;
  reg [63:0] gemm_slot_src1;
  reg [63:0] gemm_slot_dst0;
  reg [63:0] gemm_slot_dst1;
  reg [31:0] gemm_slot_size0;
  reg [31:0] gemm_slot_size1;
  reg [8:0]  gemm_slot_beats0;
  reg [8:0]  gemm_slot_beats1;
  reg [7:0]  gemm_slot_arlen0;
  reg [7:0]  gemm_slot_arlen1;
  reg        gemm_dma_sel;
  reg        gemm_done_pulse;
  reg [63:0] gemm_done_uid;
  reg [15:0] gemm_mac_a_vec0;
  reg [15:0] gemm_mac_b_vec0;
  reg [15:0] gemm_mac_a_vec1;
  reg [15:0] gemm_mac_b_vec1;
  reg signed [31:0] gemm_slot_accum0;
  reg signed [31:0] gemm_slot_accum1;
  reg [7:0] vec_in0;
  reg [7:0] vec_in1;
  reg [7:0] vec_last_result;
  reg [3:0] vec_op_sel;
  reg [3:0] vec_dtype_sel;
  reg vec_pending;
  reg vec_done_pulse;
  reg [255:0] dma_buf;
  reg [8:0]  dma_beats;
  reg [8:0]  dma_beats_left;
  reg [7:0]  dma_arlen;
  reg [255:0] dma_buf_mem [0:255];
  reg [7:0]  dma_rd_idx;
  reg [7:0]  dma_wr_idx;
  reg [31:0] error_code;

  localparam STATUS_IDLE = 32'h1;
  localparam STATUS_BUSY = 32'h2;
  localparam STATUS_ERR  = 32'h4;

  localparam integer AXI_BEAT_BYTES = 32;

  localparam IRQ_CQ_EMPTY    = 0;
  localparam IRQ_EVENT       = 1;
  localparam IRQ_ERROR       = 2;
  localparam [3:0] VEC_OP_RELU      = 4'h0;
  localparam [3:0] VEC_OP_ADD       = 4'h1;
  localparam [3:0] VEC_OP_MUL       = 4'h2;
  localparam [3:0] VEC_OP_GELU      = 4'h3;
  localparam [3:0] VEC_OP_SOFTMAX   = 4'h4;
  localparam [3:0] VEC_OP_LAYERNORM = 4'h5;
  localparam [3:0] VEC_OP_DRELU     = 4'h6;
  localparam [3:0] VEC_OP_DGELU     = 4'h7;
  localparam [3:0] VEC_OP_DSOFTMAX  = 4'h8;
  localparam [3:0] VEC_OP_DLAYERNORM= 4'h9;
  localparam [3:0] VEC_DTYPE_INT8   = 4'h0;
  localparam [3:0] VEC_DTYPE_FP16   = 4'h1;
  localparam       VEC_EN_ADD       = 1;
  localparam       VEC_EN_MUL       = 1;
  localparam       VEC_EN_RELU      = 1;
  localparam       VEC_EN_GELU      = 0;
  localparam       VEC_EN_SOFTMAX   = 0;
  localparam       VEC_EN_LAYERNORM = 0;
  localparam       VEC_EN_DRELU     = 0;
  localparam       VEC_EN_DGELU     = 0;
  localparam       VEC_EN_DSOFTMAX  = 0;
  localparam       VEC_EN_DLAYERNORM= 0;
  localparam       VEC_FP16_ENABLED = 0;
  localparam integer GEMM_MAC_LANES = 1;
  localparam integer GEMM_ELEM_BITS = 16;
  localparam integer GEMM_FP16_RAW16_PLACEHOLDER = 1;
  localparam integer GEMM_FP16_ACCUM_FP32 = 0;
  localparam integer VEC_LANES      = 1;

  // MMIO offsets (bytes)
  `include "mmio_map.vh"

  wire signed [31:0] gemm_mac_dot0;
  wire signed [31:0] gemm_mac_dot1;

  gemm_mac_fp16 #(
    .LANES(1),
    .ACC_WIDTH(32)
  ) u_gemm_mac0 (
    .a_vec(gemm_mac_a_vec0),
    .b_vec(gemm_mac_b_vec0),
    .acc_out(gemm_mac_dot0)
  );

  gemm_mac_fp16 #(
    .LANES(1),
    .ACC_WIDTH(32)
  ) u_gemm_mac1 (
    .a_vec(gemm_mac_a_vec1),
    .b_vec(gemm_mac_b_vec1),
    .acc_out(gemm_mac_dot1)
  );

  wire [7:0] vec_add_res;
  wire [7:0] vec_mul_res;
  wire [7:0] vec_relu_res;
  wire [7:0] vec_gelu_res;
  wire [7:0] vec_softmax_res;
  wire [7:0] vec_layernorm_res;
  wire [7:0] vec_drelu_res;
  wire [7:0] vec_dgelu_res;
  wire [7:0] vec_dsoftmax_res;
  wire [7:0] vec_dlayernorm_res;
  wire [7:0] vec_result_next_int8;
  wire [7:0] vec_result_next_fp16;
  wire [7:0] vec_result_next;
  wire vec_dtype_is_fp16;

  genvar gi;
  generate
    for (gi = 0; gi < 1; gi = gi + 1) begin : g_vec_lane
      assign vec_add_res[(gi*8) +: 8] = $signed(vec_in0[(gi*8) +: 8]) + $signed(vec_in1[(gi*8) +: 8]);
      assign vec_mul_res[(gi*8) +: 8] = $signed(vec_in0[(gi*8) +: 8]) * $signed(vec_in1[(gi*8) +: 8]);
      assign vec_relu_res[(gi*8) +: 8] = vec_in0[(gi*8)+7] ? 8'h00 : vec_in0[(gi*8) +: 8];
      assign vec_gelu_res[(gi*8) +: 8] = vec_in0[(gi*8)+7] ? 8'h00 : ($signed(vec_in0[(gi*8) +: 8]) >>> 1);
      assign vec_softmax_res[(gi*8) +: 8] = vec_in0[(gi*8)+7] ? 8'h00 : (($signed(vec_in0[(gi*8) +: 8]) > 8'sd31) ? 8'd127 : (vec_in0[(gi*8) +: 8] << 2));
      assign vec_layernorm_res[(gi*8) +: 8] = $signed(vec_in0[(gi*8) +: 8]) >>> 1;
      assign vec_drelu_res[(gi*8) +: 8] = ($signed(vec_in0[(gi*8) +: 8]) > 0) ? 8'h01 : 8'h00;
      assign vec_dgelu_res[(gi*8) +: 8] = ($signed(vec_in0[(gi*8) +: 8]) > 0) ? 8'h01 : 8'h00;
      wire [7:0] vec_dsoftmax_p = vec_softmax_res[(gi*8) +: 8];
      wire [15:0] vec_dsoftmax_mul = vec_dsoftmax_p * (8'd127 - vec_dsoftmax_p);
      assign vec_dsoftmax_res[(gi*8) +: 8] = vec_dsoftmax_mul[14:7];
      assign vec_dlayernorm_res[(gi*8) +: 8] = 8'h01;
    end
  endgenerate


  wire [7:0] vec_add_res_fp16 = {8{1'b0}};
  wire [7:0] vec_mul_res_fp16 = {8{1'b0}};
  wire [7:0] vec_relu_res_fp16 = {8{1'b0}};
  wire [7:0] vec_gelu_res_fp16 = {8{1'b0}};
  wire [7:0] vec_softmax_res_fp16 = {8{1'b0}};
  wire [7:0] vec_layernorm_res_fp16 = {8{1'b0}};
  wire [7:0] vec_drelu_res_fp16 = {8{1'b0}};
  wire [7:0] vec_dgelu_res_fp16 = {8{1'b0}};
  wire [7:0] vec_dsoftmax_res_fp16 = {8{1'b0}};
  wire [7:0] vec_dlayernorm_res_fp16 = {8{1'b0}};

  assign vec_dtype_is_fp16 = (vec_dtype_sel == VEC_DTYPE_FP16);

  assign vec_result_next_int8 = (vec_op_sel == VEC_OP_ADD) ? vec_add_res :
                                (vec_op_sel == VEC_OP_MUL) ? vec_mul_res :
                                (vec_op_sel == VEC_OP_GELU) ? vec_gelu_res :
                                (vec_op_sel == VEC_OP_SOFTMAX) ? vec_softmax_res :
                                (vec_op_sel == VEC_OP_LAYERNORM) ? vec_layernorm_res :
                                (vec_op_sel == VEC_OP_DRELU) ? vec_drelu_res :
                                (vec_op_sel == VEC_OP_DGELU) ? vec_dgelu_res :
                                (vec_op_sel == VEC_OP_DSOFTMAX) ? vec_dsoftmax_res :
                                (vec_op_sel == VEC_OP_DLAYERNORM) ? vec_dlayernorm_res :
                                vec_relu_res;

  assign vec_result_next_fp16 = (vec_op_sel == VEC_OP_ADD) ? vec_add_res_fp16 :
                                (vec_op_sel == VEC_OP_MUL) ? vec_mul_res_fp16 :
                                (vec_op_sel == VEC_OP_GELU) ? vec_gelu_res_fp16 :
                                (vec_op_sel == VEC_OP_SOFTMAX) ? vec_softmax_res_fp16 :
                                (vec_op_sel == VEC_OP_LAYERNORM) ? vec_layernorm_res_fp16 :
                                (vec_op_sel == VEC_OP_DRELU) ? vec_drelu_res_fp16 :
                                (vec_op_sel == VEC_OP_DGELU) ? vec_dgelu_res_fp16 :
                                (vec_op_sel == VEC_OP_DSOFTMAX) ? vec_dsoftmax_res_fp16 :
                                (vec_op_sel == VEC_OP_DLAYERNORM) ? vec_dlayernorm_res_fp16 :
                                vec_relu_res_fp16;

  assign vec_result_next = vec_dtype_is_fp16 ? vec_result_next_fp16 : vec_result_next_int8;


  always @(*) begin
    case (mmio_addr)
      OFF_VERSION:    mmio_rdata = version;
      OFF_CAPS:       mmio_rdata = capabilities;
      OFF_STATUS:     mmio_rdata = status;
      OFF_CONTROL:    mmio_rdata = control;
      OFF_IRQ_STATUS: mmio_rdata = irq_status;
      OFF_IRQ_ENABLE: mmio_rdata = irq_enable;
      OFF_CQ_BASE_LO: mmio_rdata = cq_base_lo;
      OFF_CQ_BASE_HI: mmio_rdata = cq_base_hi;
      OFF_CQ_SIZE:    mmio_rdata = cq_size;
      OFF_CQ_HEAD:    mmio_rdata = cq_head;
      OFF_CQ_TAIL:    mmio_rdata = cq_tail;
      OFF_ERROR_CODE: mmio_rdata = error_code;
      default: mmio_rdata = 0;
    endcase
  end

  always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      version <= 32'h0001_0001;
      capabilities <= 32'h0000_0133; // DMA_COPY/STRIDED/GATHER/SCATTER + GEMM/VEC/SOFTMAX + EVENT_IRQ
      status <= STATUS_IDLE;
      control <= 0;
      irq_status <= 0;
      irq_enable <= 0;
      cq_base_lo <= 0;
      cq_base_hi <= 0;
      cq_size <= 0;
      cq_head <= 0;
      cq_tail <= 0;
      cq_count <= 0;
      cq_word0 <= 0;
      cq_word0_size <= 0;
      cq_pending_ext <= 0;
      error_code <= 0;
      irq <= 0;
      last_opcode <= 0;
      last_tag <= 0;
      last_src <= 0;
      last_dst <= 0;
      last_size <= 0;
      last_op_uid <= 0;
      dma_src <= 0;
      dma_dst <= 0;
      dma_size <= 0;
      cq_stage_valid <= 0;
      dma_pending <= 0;
      dma_state <= 0;
      gemm_pending <= 0;
      gemm_slot_valid <= 0;
      gemm_slot_done <= 0;
      gemm_slot_cycles0 <= 0;
      gemm_slot_cycles1 <= 0;
      gemm_slot_uid0 <= 0;
      gemm_slot_uid1 <= 0;
      gemm_slot_src0 <= 0;
      gemm_slot_src1 <= 0;
      gemm_slot_dst0 <= 0;
      gemm_slot_dst1 <= 0;
      gemm_slot_size0 <= 0;
      gemm_slot_size1 <= 0;
      gemm_slot_beats0 <= 0;
      gemm_slot_beats1 <= 0;
      gemm_slot_arlen0 <= 0;
      gemm_slot_arlen1 <= 0;
      gemm_dma_sel <= 0;
      gemm_done_pulse <= 0;
      gemm_done_uid <= 0;
      gemm_mac_a_vec0 <= 0;
      gemm_mac_b_vec0 <= 0;
      gemm_mac_a_vec1 <= 0;
      gemm_mac_b_vec1 <= 0;
      gemm_slot_accum0 <= 0;
      gemm_slot_accum1 <= 0;
      vec_in0 <= 0;
      vec_in1 <= 0;
      vec_last_result <= 0;
      vec_op_sel <= 0;
      vec_dtype_sel <= 0;
      vec_pending <= 0;
      vec_done_pulse <= 0;
      dma_buf <= 0;
      dma_beats <= 0;
      dma_beats_left <= 0;
      dma_arlen <= 0;
      dma_rd_idx <= 0;
      dma_wr_idx <= 0;
      dma_req_valid <= 0;
      dma_req_src <= 0;
      dma_req_dst <= 0;
      dma_req_bytes <= 0;
      m_axi_awvalid <= 1'b0;
      m_axi_awaddr <= 0;
      m_axi_awlen <= 0;
      m_axi_awsize <= 0;
      m_axi_wvalid <= 1'b0;
      m_axi_wdata <= 0;
      m_axi_wstrb <= 0;
      m_axi_wlast <= 1'b0;
      m_axi_bready <= 1'b0;
      m_axi_arvalid <= 1'b0;
      m_axi_araddr <= 0;
      m_axi_arlen <= 0;
      m_axi_arsize <= 0;
      m_axi_rready <= 1'b0;
    end else begin
      // Default: clear level IRQ unless status bit set
      irq <= |(irq_status & irq_enable);
      if (dma_req_valid && dma_req_ready) begin
        dma_req_valid <= 0;
      end
      if (dma_resp_done) begin
        irq_status[IRQ_EVENT] <= 1'b1;
      end
      // Two-slot GEMM stub with OOO-capable completion scheduling.
      gemm_done_pulse <= 1'b0;
      vec_done_pulse <= 1'b0;
      if (vec_pending) begin
        vec_last_result <= vec_result_next;
        vec_pending <= 1'b0;
        vec_done_pulse <= 1'b1;
        irq_status[IRQ_EVENT] <= 1'b1;
      end
      if (gemm_slot_valid[0] && !gemm_slot_done[0]) begin
        gemm_slot_accum0 <= gemm_slot_accum0 + gemm_mac_dot0;
      end
      if (gemm_slot_valid[1] && !gemm_slot_done[1]) begin
        gemm_slot_accum1 <= gemm_slot_accum1 + gemm_mac_dot1;
      end
      if (gemm_slot_valid[0] && !gemm_slot_done[0]) begin
        if (gemm_slot_cycles0 != 0) begin
          gemm_slot_cycles0 <= gemm_slot_cycles0 - 1;
          if (gemm_slot_cycles0 == 1) begin
            gemm_slot_done[0] <= 1'b1;
            gemm_done_pulse <= 1'b1;
            gemm_done_uid <= gemm_slot_uid0;
          end
        end else begin
          gemm_slot_done[0] <= 1'b1;
          gemm_done_pulse <= 1'b1;
          gemm_done_uid <= gemm_slot_uid0;
        end
      end
      if (gemm_slot_valid[1] && !gemm_slot_done[1]) begin
        if (gemm_slot_cycles1 != 0) begin
          gemm_slot_cycles1 <= gemm_slot_cycles1 - 1;
          if (gemm_slot_cycles1 == 1) begin
            gemm_slot_done[1] <= 1'b1;
            gemm_done_pulse <= 1'b1;
            gemm_done_uid <= gemm_slot_uid1;
          end
        end else begin
          gemm_slot_done[1] <= 1'b1;
          gemm_done_pulse <= 1'b1;
          gemm_done_uid <= gemm_slot_uid1;
        end
      end
      // Prefer slot1 if both are done, so completion order can differ from issue order.
      if (!dma_pending) begin
        if (gemm_slot_done[1]) begin
          dma_src <= gemm_slot_src1;
          dma_dst <= gemm_slot_dst1;
          dma_size <= gemm_slot_size1;
          dma_beats <= gemm_slot_beats1;
          dma_arlen <= gemm_slot_arlen1;
          dma_pending <= 1'b1;
          gemm_slot_valid[1] <= 1'b0;
          gemm_slot_done[1] <= 1'b0;
          gemm_dma_sel <= 1'b1;
        end else if (gemm_slot_done[0]) begin
          dma_src <= gemm_slot_src0;
          dma_dst <= gemm_slot_dst0;
          dma_size <= gemm_slot_size0;
          dma_beats <= gemm_slot_beats0;
          dma_arlen <= gemm_slot_arlen0;
          dma_pending <= 1'b1;
          gemm_slot_valid[0] <= 1'b0;
          gemm_slot_done[0] <= 1'b0;
          gemm_dma_sel <= 1'b0;
        end
      end
      gemm_pending <= (gemm_slot_valid != 2'b00);
      m_axi_awvalid <= 1'b0;
      m_axi_awaddr <= 0;
      m_axi_awlen <= 0;
      m_axi_awsize <= 0;
      m_axi_wvalid <= 1'b0;
      m_axi_wdata <= 0;
      m_axi_wstrb <= 0;
      m_axi_wlast <= 1'b0;
      m_axi_bready <= 1'b0;
      m_axi_arvalid <= 1'b0;
      m_axi_araddr <= 0;
      m_axi_arlen <= 0;
      m_axi_arsize <= 0;
      m_axi_rready <= 1'b0;
      // AXI DMA shim: burst read then burst write.
      case (dma_state)
        0: begin
          if (dma_pending) begin
            if (dma_beats_left == 0) begin
              dma_beats_left <= dma_beats;
              dma_rd_idx <= 0;
              dma_wr_idx <= 0;
            end
            m_axi_arvalid <= 1'b1;
            m_axi_araddr <= dma_src;
            m_axi_arlen <= dma_arlen;
            m_axi_arsize <= 3'd5; // beat bytes = 2**5
            if (m_axi_arready) begin
              dma_state <= 1;
            end
          end
        end
        1: begin
          m_axi_rready <= 1'b1;
          if (m_axi_rvalid) begin
            dma_buf_mem[dma_rd_idx] <= m_axi_rdata;
            dma_rd_idx <= dma_rd_idx + 1;
            if (m_axi_rlast) begin
              dma_state <= 2;
            end
          end
        end
        2: begin
          m_axi_awvalid <= 1'b1;
          m_axi_awaddr <= dma_dst;
          m_axi_awlen <= dma_arlen;
          m_axi_awsize <= 3'd5;
          if (m_axi_awready) begin
            dma_state <= 3;
          end
        end
        3: begin
          m_axi_wvalid <= 1'b1;
          m_axi_wdata <= dma_buf_mem[dma_wr_idx];
          m_axi_wstrb <= {32{1'b1}};
          m_axi_wlast <= (dma_beats_left == 1);
          if (m_axi_wready) begin
            if (dma_beats_left == 1) begin
              dma_state <= 4;
            end else begin
              dma_wr_idx <= dma_wr_idx + 1;
              dma_beats_left <= dma_beats_left - 1;
            end
          end
        end
        4: begin
          m_axi_bready <= 1'b1;
          if (m_axi_bvalid) begin
            dma_beats_left <= 0;
            dma_state <= 0;
            dma_pending <= 1'b0;
            irq_status[IRQ_EVENT] <= 1'b1;
          end
        end
        default: dma_state <= 0;
      endcase

      if (mmio_we) begin
        case (mmio_addr)
          OFF_CONTROL: control <= mmio_wdata;
          OFF_IRQ_STATUS: irq_status <= irq_status & ~mmio_wdata; // W1C
          OFF_IRQ_ENABLE: irq_enable <= mmio_wdata;
          OFF_CQ_BASE_LO: cq_base_lo <= mmio_wdata;
          OFF_CQ_BASE_HI: cq_base_hi <= mmio_wdata;
          OFF_CQ_SIZE:    cq_size <= mmio_wdata;
          OFF_CQ_TAIL:    cq_tail <= mmio_wdata;
          OFF_DOORBELL: begin
            // Minimal behavior: consume all queued descriptors.
            cq_count <= ((cq_tail - cq_head) >> 5);
            if (((cq_tail - cq_head) >> 5) == 0) begin
              status <= STATUS_IDLE;
              irq_status[IRQ_CQ_EMPTY] <= 1'b1;
            end else begin
              status <= STATUS_BUSY;
            end
            // DMA request will be issued when DMA_COPY descriptor is fetched.
          end
          default: begin end
        endcase
      end

      // Command queue fetch (supports v0.1 32B and v0.2 64B descriptors).
      if (cq_count != 0) begin
        if (!cq_stage_valid && !cq_pending_ext) begin
          cq_mem_addr <= {cq_base_hi, cq_base_lo} + cq_head;
          cq_stage_valid <= 1'b1;
        end else if (cq_stage_valid && !cq_pending_ext) begin
          cq_word0 <= cq_mem_rdata;
          cq_word0_size <= cq_mem_rdata[23:16];
          if (cq_mem_rdata[23:16] >= 8'h02) begin
            cq_pending_ext <= 1'b1;
            cq_stage_valid <= 1'b0;
          end else begin
            last_opcode <= cq_mem_rdata[7:0];
            last_tag <= cq_mem_rdata[63:32];
            last_src <= cq_mem_rdata[127:64];
            last_dst <= cq_mem_rdata[191:128];
            last_size <= cq_mem_rdata[223:192];
            last_op_uid <= 0;
            if (cq_mem_rdata[7:0] == 8'h01) begin
              dma_req_valid <= 1'b1;
              dma_req_src <= cq_mem_rdata[127:64];
              dma_req_dst <= cq_mem_rdata[191:128];
              dma_req_bytes <= cq_mem_rdata[223:192];
              dma_src <= cq_mem_rdata[127:64];
              dma_dst <= cq_mem_rdata[191:128];
              dma_size <= cq_mem_rdata[223:192];
              dma_beats <= (cq_mem_rdata[223:197] + (|cq_mem_rdata[196:192]));
              dma_arlen <= (cq_mem_rdata[223:197] + (|cq_mem_rdata[196:192])) - 1;
              dma_pending <= 1'b1;
            end else if (cq_mem_rdata[7:0] == 8'h10) begin
              // GEMM stub: v0.1 sizes packed in TAG.
              if (!gemm_slot_valid[0]) begin
                gemm_slot_valid[0] <= 1'b1;
                gemm_slot_done[0] <= 1'b0;
                gemm_slot_uid0 <= 64'h0;
                gemm_mac_a_vec0 <= cq_mem_rdata[79:64];
                gemm_mac_b_vec0 <= cq_mem_rdata[143:128];
                gemm_slot_accum0 <= 0;
                if ((cq_mem_rdata[63:52] == 0) || (cq_mem_rdata[51:42] == 0) || (cq_mem_rdata[41:32] == 0)) begin
                  gemm_slot_cycles0 <= 1;
                end else begin
                  gemm_slot_cycles0 <= (((cq_mem_rdata[63:52] * cq_mem_rdata[51:42] * cq_mem_rdata[41:32]) >> 10) + 1);
                end
                gemm_slot_src0 <= cq_mem_rdata[127:64];
                gemm_slot_dst0 <= cq_mem_rdata[255:192];
                gemm_slot_size0 <= ((cq_mem_rdata[11:8] == 4'h1 || cq_mem_rdata[11:8] == 4'h2)
                                    ? (cq_mem_rdata[63:52] * cq_mem_rdata[51:42] * 2)
                                    : (cq_mem_rdata[63:52] * cq_mem_rdata[51:42]));
                gemm_slot_beats0 <= (((((cq_mem_rdata[11:8] == 4'h1 || cq_mem_rdata[11:8] == 4'h2)
                                        ? (cq_mem_rdata[63:52] * cq_mem_rdata[51:42] * 2)
                                        : (cq_mem_rdata[63:52] * cq_mem_rdata[51:42]))
                                       + AXI_BEAT_BYTES - 1) >> 5));
                gemm_slot_arlen0 <= (((((cq_mem_rdata[11:8] == 4'h1 || cq_mem_rdata[11:8] == 4'h2)
                                        ? (cq_mem_rdata[63:52] * cq_mem_rdata[51:42] * 2)
                                        : (cq_mem_rdata[63:52] * cq_mem_rdata[51:42]))
                                       + AXI_BEAT_BYTES - 1) >> 5) - 1);
              end else if (!gemm_slot_valid[1]) begin
                gemm_slot_valid[1] <= 1'b1;
                gemm_slot_done[1] <= 1'b0;
                gemm_slot_uid1 <= 64'h0;
                gemm_mac_a_vec1 <= cq_mem_rdata[79:64];
                gemm_mac_b_vec1 <= cq_mem_rdata[143:128];
                gemm_slot_accum1 <= 0;
                if ((cq_mem_rdata[63:52] == 0) || (cq_mem_rdata[51:42] == 0) || (cq_mem_rdata[41:32] == 0)) begin
                  gemm_slot_cycles1 <= 1;
                end else begin
                  gemm_slot_cycles1 <= (((cq_mem_rdata[63:52] * cq_mem_rdata[51:42] * cq_mem_rdata[41:32]) >> 10) + 1);
                end
                gemm_slot_src1 <= cq_mem_rdata[127:64];
                gemm_slot_dst1 <= cq_mem_rdata[255:192];
                gemm_slot_size1 <= ((cq_mem_rdata[11:8] == 4'h1 || cq_mem_rdata[11:8] == 4'h2)
                                    ? (cq_mem_rdata[63:52] * cq_mem_rdata[51:42] * 2)
                                    : (cq_mem_rdata[63:52] * cq_mem_rdata[51:42]));
                gemm_slot_beats1 <= (((((cq_mem_rdata[11:8] == 4'h1 || cq_mem_rdata[11:8] == 4'h2)
                                        ? (cq_mem_rdata[63:52] * cq_mem_rdata[51:42] * 2)
                                        : (cq_mem_rdata[63:52] * cq_mem_rdata[51:42]))
                                       + AXI_BEAT_BYTES - 1) >> 5));
                gemm_slot_arlen1 <= (((((cq_mem_rdata[11:8] == 4'h1 || cq_mem_rdata[11:8] == 4'h2)
                                        ? (cq_mem_rdata[63:52] * cq_mem_rdata[51:42] * 2)
                                        : (cq_mem_rdata[63:52] * cq_mem_rdata[51:42]))
                                       + AXI_BEAT_BYTES - 1) >> 5) - 1);
              end else begin
                error_code <= 32'h2; // GEMM in-flight queue full
              end
            end else if (cq_mem_rdata[7:0] == 8'h11) begin
              // VEC_OP (v0.1): input vectors are carried in descriptor payload bytes.
              if (vec_pending) begin
                error_code <= 32'h3; // VEC in-flight queue full
              end else begin
                vec_in0 <= cq_mem_rdata[71:64];
                vec_in1 <= cq_mem_rdata[135:128];
                vec_op_sel <= cq_mem_rdata[11:8];
                vec_dtype_sel <= cq_mem_rdata[15:12];
                if (((cq_mem_rdata[15:12] == VEC_DTYPE_FP16) && !VEC_FP16_ENABLED) ||
                    ((cq_mem_rdata[15:12] != VEC_DTYPE_INT8) && (cq_mem_rdata[15:12] != VEC_DTYPE_FP16)) ||
                    ((cq_mem_rdata[15:12] == VEC_DTYPE_FP16) &&
                     (cq_mem_rdata[11:8] != VEC_OP_RELU) &&
                     (cq_mem_rdata[11:8] != VEC_OP_ADD) &&
                     (cq_mem_rdata[11:8] != VEC_OP_MUL) &&
                     (cq_mem_rdata[11:8] != VEC_OP_GELU) &&
                     (cq_mem_rdata[11:8] != VEC_OP_SOFTMAX) &&
                     (cq_mem_rdata[11:8] != VEC_OP_LAYERNORM) &&
                     (cq_mem_rdata[11:8] != VEC_OP_DRELU) &&
                     (cq_mem_rdata[11:8] != VEC_OP_DGELU) &&
                     (cq_mem_rdata[11:8] != VEC_OP_DSOFTMAX) &&
                     (cq_mem_rdata[11:8] != VEC_OP_DLAYERNORM)) ||
                    (cq_mem_rdata[11:8] == VEC_OP_ADD       && !VEC_EN_ADD)       ||
                    (cq_mem_rdata[11:8] == VEC_OP_MUL       && !VEC_EN_MUL)       ||
                    (cq_mem_rdata[11:8] == VEC_OP_RELU      && !VEC_EN_RELU)      ||
                    (cq_mem_rdata[11:8] == VEC_OP_GELU      && !VEC_EN_GELU)      ||
                    (cq_mem_rdata[11:8] == VEC_OP_SOFTMAX   && !VEC_EN_SOFTMAX)   ||
                    (cq_mem_rdata[11:8] == VEC_OP_LAYERNORM && !VEC_EN_LAYERNORM) ||
                    (cq_mem_rdata[11:8] == VEC_OP_DRELU     && !VEC_EN_DRELU)     ||
                    (cq_mem_rdata[11:8] == VEC_OP_DGELU     && !VEC_EN_DGELU)     ||
                    (cq_mem_rdata[11:8] == VEC_OP_DSOFTMAX  && !VEC_EN_DSOFTMAX)  ||
                    (cq_mem_rdata[11:8] == VEC_OP_DLAYERNORM&& !VEC_EN_DLAYERNORM)||
                    ((cq_mem_rdata[11:8] != VEC_OP_RELU)      &&
                     (cq_mem_rdata[11:8] != VEC_OP_ADD)       &&
                     (cq_mem_rdata[11:8] != VEC_OP_MUL)       &&
                     (cq_mem_rdata[11:8] != VEC_OP_GELU)      &&
                     (cq_mem_rdata[11:8] != VEC_OP_SOFTMAX)   &&
                     (cq_mem_rdata[11:8] != VEC_OP_LAYERNORM) &&
                     (cq_mem_rdata[11:8] != VEC_OP_DRELU)     &&
                     (cq_mem_rdata[11:8] != VEC_OP_DGELU)     &&
                     (cq_mem_rdata[11:8] != VEC_OP_DSOFTMAX)  &&
                     (cq_mem_rdata[11:8] != VEC_OP_DLAYERNORM))) begin
                  error_code <= 32'h6; // unsupported configured VEC op
                end else begin
                  vec_pending <= 1'b1;
                end
              end
            end else if (cq_mem_rdata[7:0] == 8'h20) begin
              // EVENT_SIGNAL: immediately signal
              irq_status[IRQ_EVENT] <= 1'b1;
            end else if (cq_mem_rdata[7:0] == 8'h21) begin
              // EVENT_WAIT: stubbed as immediately satisfied
              irq_status[IRQ_EVENT] <= 1'b1;
            end else begin
              error_code <= 32'h1;
            end
            cq_head <= cq_head + 32;
            if (cq_count == 1) begin
              irq_status[IRQ_CQ_EMPTY] <= 1'b1;
            end
            cq_count <= cq_count - 1;
            cq_stage_valid <= 1'b0;
          end
        end else if (cq_pending_ext) begin
          if (!cq_stage_valid) begin
            cq_mem_addr <= {cq_base_hi, cq_base_lo} + cq_head + 32;
            cq_stage_valid <= 1'b1;
          end else begin
            last_opcode <= cq_word0[7:0];
            last_tag <= cq_word0[63:32];
            last_src <= cq_word0[127:64];
            last_dst <= cq_word0[191:128];
            last_size <= cq_mem_rdata[31:0];
            last_op_uid <= cq_mem_rdata[255:192];
            if (cq_word0[7:0] == 8'h10) begin
              // GEMM stub: v0.2 sizes in extension.
              if (!gemm_slot_valid[0]) begin
                gemm_slot_valid[0] <= 1'b1;
                gemm_slot_done[0] <= 1'b0;
                gemm_slot_uid0 <= cq_mem_rdata[255:192];
                gemm_mac_a_vec0 <= cq_word0[79:64];
                gemm_mac_b_vec0 <= cq_word0[143:128];
                gemm_slot_accum0 <= 0;
                if ((cq_mem_rdata[31:0] == 0) || (cq_mem_rdata[63:32] == 0) || (cq_mem_rdata[95:64] == 0)) begin
                  gemm_slot_cycles0 <= 1;
                end else begin
                  // Optional UID-based jitter (bit63) to exercise OOO completion in tests.
                  gemm_slot_cycles0 <= (((cq_mem_rdata[31:0] * cq_mem_rdata[63:32] * cq_mem_rdata[95:64]) >> 10)
                                        + 1 + (cq_mem_rdata[255] ? 8 : 0));
                end
                gemm_slot_src0 <= cq_word0[127:64];
                gemm_slot_dst0 <= cq_word0[255:192];
                gemm_slot_size0 <= ((cq_word0[11:8] == 4'h1 || cq_word0[11:8] == 4'h2)
                                    ? (cq_mem_rdata[31:0] * cq_mem_rdata[63:32] * 2)
                                    : (cq_mem_rdata[31:0] * cq_mem_rdata[63:32]));
                gemm_slot_beats0 <= (((((cq_word0[11:8] == 4'h1 || cq_word0[11:8] == 4'h2)
                                        ? (cq_mem_rdata[31:0] * cq_mem_rdata[63:32] * 2)
                                        : (cq_mem_rdata[31:0] * cq_mem_rdata[63:32]))
                                       + AXI_BEAT_BYTES - 1) >> 5));
                gemm_slot_arlen0 <= (((((cq_word0[11:8] == 4'h1 || cq_word0[11:8] == 4'h2)
                                        ? (cq_mem_rdata[31:0] * cq_mem_rdata[63:32] * 2)
                                        : (cq_mem_rdata[31:0] * cq_mem_rdata[63:32]))
                                       + AXI_BEAT_BYTES - 1) >> 5) - 1);
              end else if (!gemm_slot_valid[1]) begin
                gemm_slot_valid[1] <= 1'b1;
                gemm_slot_done[1] <= 1'b0;
                gemm_slot_uid1 <= cq_mem_rdata[255:192];
                gemm_mac_a_vec1 <= cq_word0[79:64];
                gemm_mac_b_vec1 <= cq_word0[143:128];
                gemm_slot_accum1 <= 0;
                if ((cq_mem_rdata[31:0] == 0) || (cq_mem_rdata[63:32] == 0) || (cq_mem_rdata[95:64] == 0)) begin
                  gemm_slot_cycles1 <= 1;
                end else begin
                  gemm_slot_cycles1 <= (((cq_mem_rdata[31:0] * cq_mem_rdata[63:32] * cq_mem_rdata[95:64]) >> 10)
                                        + 1 + (cq_mem_rdata[255] ? 8 : 0));
                end
                gemm_slot_src1 <= cq_word0[127:64];
                gemm_slot_dst1 <= cq_word0[255:192];
                gemm_slot_size1 <= ((cq_word0[11:8] == 4'h1 || cq_word0[11:8] == 4'h2)
                                    ? (cq_mem_rdata[31:0] * cq_mem_rdata[63:32] * 2)
                                    : (cq_mem_rdata[31:0] * cq_mem_rdata[63:32]));
                gemm_slot_beats1 <= (((((cq_word0[11:8] == 4'h1 || cq_word0[11:8] == 4'h2)
                                        ? (cq_mem_rdata[31:0] * cq_mem_rdata[63:32] * 2)
                                        : (cq_mem_rdata[31:0] * cq_mem_rdata[63:32]))
                                       + AXI_BEAT_BYTES - 1) >> 5));
                gemm_slot_arlen1 <= (((((cq_word0[11:8] == 4'h1 || cq_word0[11:8] == 4'h2)
                                        ? (cq_mem_rdata[31:0] * cq_mem_rdata[63:32] * 2)
                                        : (cq_mem_rdata[31:0] * cq_mem_rdata[63:32]))
                                       + AXI_BEAT_BYTES - 1) >> 5) - 1);
              end else begin
                error_code <= 32'h2; // GEMM in-flight queue full
              end
            end else if (cq_word0[7:0] == 8'h11) begin
              // VEC_OP (v0.2 base word): vectors are sourced from header payload.
              if (vec_pending) begin
                error_code <= 32'h3; // VEC in-flight queue full
              end else begin
                vec_in0 <= cq_word0[71:64];
                vec_in1 <= cq_word0[135:128];
                vec_op_sel <= cq_word0[11:8];
                vec_dtype_sel <= cq_word0[15:12];
                if (((cq_word0[15:12] == VEC_DTYPE_FP16) && !VEC_FP16_ENABLED) ||
                    ((cq_word0[15:12] != VEC_DTYPE_INT8) && (cq_word0[15:12] != VEC_DTYPE_FP16)) ||
                    ((cq_word0[15:12] == VEC_DTYPE_FP16) &&
                     (cq_word0[11:8] != VEC_OP_RELU) &&
                     (cq_word0[11:8] != VEC_OP_ADD) &&
                     (cq_word0[11:8] != VEC_OP_MUL) &&
                     (cq_word0[11:8] != VEC_OP_GELU) &&
                     (cq_word0[11:8] != VEC_OP_SOFTMAX) &&
                     (cq_word0[11:8] != VEC_OP_LAYERNORM) &&
                     (cq_word0[11:8] != VEC_OP_DRELU) &&
                     (cq_word0[11:8] != VEC_OP_DGELU) &&
                     (cq_word0[11:8] != VEC_OP_DSOFTMAX) &&
                     (cq_word0[11:8] != VEC_OP_DLAYERNORM)) ||
                    (cq_word0[11:8] == VEC_OP_ADD       && !VEC_EN_ADD)       ||
                    (cq_word0[11:8] == VEC_OP_MUL       && !VEC_EN_MUL)       ||
                    (cq_word0[11:8] == VEC_OP_RELU      && !VEC_EN_RELU)      ||
                    (cq_word0[11:8] == VEC_OP_GELU      && !VEC_EN_GELU)      ||
                    (cq_word0[11:8] == VEC_OP_SOFTMAX   && !VEC_EN_SOFTMAX)   ||
                    (cq_word0[11:8] == VEC_OP_LAYERNORM && !VEC_EN_LAYERNORM) ||
                    (cq_word0[11:8] == VEC_OP_DRELU     && !VEC_EN_DRELU)     ||
                    (cq_word0[11:8] == VEC_OP_DGELU     && !VEC_EN_DGELU)     ||
                    (cq_word0[11:8] == VEC_OP_DSOFTMAX  && !VEC_EN_DSOFTMAX)  ||
                    (cq_word0[11:8] == VEC_OP_DLAYERNORM&& !VEC_EN_DLAYERNORM)||
                    ((cq_word0[11:8] != VEC_OP_RELU)      &&
                     (cq_word0[11:8] != VEC_OP_ADD)       &&
                     (cq_word0[11:8] != VEC_OP_MUL)       &&
                     (cq_word0[11:8] != VEC_OP_GELU)      &&
                     (cq_word0[11:8] != VEC_OP_SOFTMAX)   &&
                     (cq_word0[11:8] != VEC_OP_LAYERNORM) &&
                     (cq_word0[11:8] != VEC_OP_DRELU)     &&
                     (cq_word0[11:8] != VEC_OP_DGELU)     &&
                     (cq_word0[11:8] != VEC_OP_DSOFTMAX)  &&
                     (cq_word0[11:8] != VEC_OP_DLAYERNORM))) begin
                  error_code <= 32'h6;
                end else begin
                  vec_pending <= 1'b1;
                end
              end
            end else begin
              error_code <= 32'h1;
            end
            if (cq_count <= cq_word0_size) begin
              irq_status[IRQ_CQ_EMPTY] <= 1'b1;
            end
            cq_head <= cq_head + (cq_word0_size * 32);
            cq_count <= cq_count - cq_word0_size;
            cq_stage_valid <= 1'b0;
            cq_pending_ext <= 1'b0;
          end
        end
      end

      if (error_code != 0) begin
        status <= STATUS_ERR;
        irq_status[IRQ_ERROR] <= 1'b1;
      end else if (!(mmio_we && mmio_addr == OFF_DOORBELL)) begin
        if ((cq_count != 0) || cq_stage_valid || dma_pending || vec_pending || (gemm_slot_valid != 2'b00)) begin
          status <= STATUS_BUSY;
        end else begin
          status <= STATUS_IDLE;
        end
      end
    end
  end

endmodule
