localparam int SRAM_COUNT = 1;
localparam int SRAM_MAX = 8;
localparam logic [63:0] SRAM_BASE0 = 64'h0000000080000000;
localparam logic [63:0] SRAM_SIZE0 = 4194304;
localparam int SRAM_ALIGN0 = 64;
localparam int SRAM_WORD_BYTES0 = 32;
localparam logic [63:0] SRAM_BASE1 = 64'h0;
localparam logic [63:0] SRAM_SIZE1 = 0;
localparam int SRAM_ALIGN1 = 0;
localparam int SRAM_WORD_BYTES1 = 0;
localparam logic [63:0] SRAM_BASE2 = 64'h0;
localparam logic [63:0] SRAM_SIZE2 = 0;
localparam int SRAM_ALIGN2 = 0;
localparam int SRAM_WORD_BYTES2 = 0;
localparam logic [63:0] SRAM_BASE3 = 64'h0;
localparam logic [63:0] SRAM_SIZE3 = 0;
localparam int SRAM_ALIGN3 = 0;
localparam int SRAM_WORD_BYTES3 = 0;
localparam logic [63:0] SRAM_BASE4 = 64'h0;
localparam logic [63:0] SRAM_SIZE4 = 0;
localparam int SRAM_ALIGN4 = 0;
localparam int SRAM_WORD_BYTES4 = 0;
localparam logic [63:0] SRAM_BASE5 = 64'h0;
localparam logic [63:0] SRAM_SIZE5 = 0;
localparam int SRAM_ALIGN5 = 0;
localparam int SRAM_WORD_BYTES5 = 0;
localparam logic [63:0] SRAM_BASE6 = 64'h0;
localparam logic [63:0] SRAM_SIZE6 = 0;
localparam int SRAM_ALIGN6 = 0;
localparam int SRAM_WORD_BYTES6 = 0;
localparam logic [63:0] SRAM_BASE7 = 64'h0;
localparam logic [63:0] SRAM_SIZE7 = 0;
localparam int SRAM_ALIGN7 = 0;
localparam int SRAM_WORD_BYTES7 = 0;
