module adder_koggestone_16u(
  input [15:0] a,
  input [15:0] b,
  output [15:0] sum,
  output cout
);

  wire p_0_0;
  wire g_0_0;
 assign p_0_0 = a[0] ^ b[0];
 assign g_0_0 = a[0] & b[0];
  wire p_1_1;
  wire g_1_1;
 assign p_1_1 = a[1] ^ b[1];
 assign g_1_1 = a[1] & b[1];
  wire p_1_0;
  wire g_1_0;
  wire p_2_2;
  wire g_2_2;
 assign p_2_2 = a[2] ^ b[2];
 assign g_2_2 = a[2] & b[2];
  wire p_2_0;
  wire g_2_0;
  wire p_2_1;
  wire g_2_1;
  wire p_3_3;
  wire g_3_3;
 assign p_3_3 = a[3] ^ b[3];
 assign g_3_3 = a[3] & b[3];
  wire p_3_0;
  wire g_3_0;
  wire p_3_1;
  wire g_3_1;
  wire p_3_2;
  wire g_3_2;
  wire p_4_4;
  wire g_4_4;
 assign p_4_4 = a[4] ^ b[4];
 assign g_4_4 = a[4] & b[4];
  wire p_4_0;
  wire g_4_0;
  wire p_4_1;
  wire g_4_1;
  wire p_4_2;
  wire g_4_2;
  wire p_4_3;
  wire g_4_3;
  wire p_5_5;
  wire g_5_5;
 assign p_5_5 = a[5] ^ b[5];
 assign g_5_5 = a[5] & b[5];
  wire p_5_0;
  wire g_5_0;
  wire p_5_1;
  wire g_5_1;
  wire p_5_2;
  wire g_5_2;
  wire p_5_3;
  wire g_5_3;
  wire p_5_4;
  wire g_5_4;
  wire p_6_6;
  wire g_6_6;
 assign p_6_6 = a[6] ^ b[6];
 assign g_6_6 = a[6] & b[6];
  wire p_6_0;
  wire g_6_0;
  wire p_6_1;
  wire g_6_1;
  wire p_6_2;
  wire g_6_2;
  wire p_6_3;
  wire g_6_3;
  wire p_6_4;
  wire g_6_4;
  wire p_6_5;
  wire g_6_5;
  wire p_7_7;
  wire g_7_7;
 assign p_7_7 = a[7] ^ b[7];
 assign g_7_7 = a[7] & b[7];
  wire p_7_0;
  wire g_7_0;
  wire p_7_1;
  wire g_7_1;
  wire p_7_2;
  wire g_7_2;
  wire p_7_3;
  wire g_7_3;
  wire p_7_4;
  wire g_7_4;
  wire p_7_5;
  wire g_7_5;
  wire p_7_6;
  wire g_7_6;
  wire p_8_8;
  wire g_8_8;
 assign p_8_8 = a[8] ^ b[8];
 assign g_8_8 = a[8] & b[8];
  wire p_8_0;
  wire g_8_0;
  wire p_8_1;
  wire g_8_1;
  wire p_8_2;
  wire g_8_2;
  wire p_8_3;
  wire g_8_3;
  wire p_8_4;
  wire g_8_4;
  wire p_8_5;
  wire g_8_5;
  wire p_8_6;
  wire g_8_6;
  wire p_8_7;
  wire g_8_7;
  wire p_9_9;
  wire g_9_9;
 assign p_9_9 = a[9] ^ b[9];
 assign g_9_9 = a[9] & b[9];
  wire p_9_0;
  wire g_9_0;
  wire p_9_1;
  wire g_9_1;
  wire p_9_2;
  wire g_9_2;
  wire p_9_3;
  wire g_9_3;
  wire p_9_4;
  wire g_9_4;
  wire p_9_5;
  wire g_9_5;
  wire p_9_6;
  wire g_9_6;
  wire p_9_7;
  wire g_9_7;
  wire p_9_8;
  wire g_9_8;
  wire p_10_10;
  wire g_10_10;
 assign p_10_10 = a[10] ^ b[10];
 assign g_10_10 = a[10] & b[10];
  wire p_10_0;
  wire g_10_0;
  wire p_10_1;
  wire g_10_1;
  wire p_10_2;
  wire g_10_2;
  wire p_10_3;
  wire g_10_3;
  wire p_10_4;
  wire g_10_4;
  wire p_10_5;
  wire g_10_5;
  wire p_10_6;
  wire g_10_6;
  wire p_10_7;
  wire g_10_7;
  wire p_10_8;
  wire g_10_8;
  wire p_10_9;
  wire g_10_9;
  wire p_11_11;
  wire g_11_11;
 assign p_11_11 = a[11] ^ b[11];
 assign g_11_11 = a[11] & b[11];
  wire p_11_0;
  wire g_11_0;
  wire p_11_1;
  wire g_11_1;
  wire p_11_2;
  wire g_11_2;
  wire p_11_3;
  wire g_11_3;
  wire p_11_4;
  wire g_11_4;
  wire p_11_5;
  wire g_11_5;
  wire p_11_6;
  wire g_11_6;
  wire p_11_7;
  wire g_11_7;
  wire p_11_8;
  wire g_11_8;
  wire p_11_9;
  wire g_11_9;
  wire p_11_10;
  wire g_11_10;
  wire p_12_12;
  wire g_12_12;
 assign p_12_12 = a[12] ^ b[12];
 assign g_12_12 = a[12] & b[12];
  wire p_12_0;
  wire g_12_0;
  wire p_12_1;
  wire g_12_1;
  wire p_12_2;
  wire g_12_2;
  wire p_12_3;
  wire g_12_3;
  wire p_12_4;
  wire g_12_4;
  wire p_12_5;
  wire g_12_5;
  wire p_12_6;
  wire g_12_6;
  wire p_12_7;
  wire g_12_7;
  wire p_12_8;
  wire g_12_8;
  wire p_12_9;
  wire g_12_9;
  wire p_12_10;
  wire g_12_10;
  wire p_12_11;
  wire g_12_11;
  wire p_13_13;
  wire g_13_13;
 assign p_13_13 = a[13] ^ b[13];
 assign g_13_13 = a[13] & b[13];
  wire p_13_0;
  wire g_13_0;
  wire p_13_1;
  wire g_13_1;
  wire p_13_2;
  wire g_13_2;
  wire p_13_3;
  wire g_13_3;
  wire p_13_4;
  wire g_13_4;
  wire p_13_5;
  wire g_13_5;
  wire p_13_6;
  wire g_13_6;
  wire p_13_7;
  wire g_13_7;
  wire p_13_8;
  wire g_13_8;
  wire p_13_9;
  wire g_13_9;
  wire p_13_10;
  wire g_13_10;
  wire p_13_11;
  wire g_13_11;
  wire p_13_12;
  wire g_13_12;
  wire p_14_14;
  wire g_14_14;
 assign p_14_14 = a[14] ^ b[14];
 assign g_14_14 = a[14] & b[14];
  wire p_14_0;
  wire g_14_0;
  wire p_14_1;
  wire g_14_1;
  wire p_14_2;
  wire g_14_2;
  wire p_14_3;
  wire g_14_3;
  wire p_14_4;
  wire g_14_4;
  wire p_14_5;
  wire g_14_5;
  wire p_14_6;
  wire g_14_6;
  wire p_14_7;
  wire g_14_7;
  wire p_14_8;
  wire g_14_8;
  wire p_14_9;
  wire g_14_9;
  wire p_14_10;
  wire g_14_10;
  wire p_14_11;
  wire g_14_11;
  wire p_14_12;
  wire g_14_12;
  wire p_14_13;
  wire g_14_13;
  wire p_15_15;
  wire g_15_15;
 assign p_15_15 = a[15] ^ b[15];
 assign g_15_15 = a[15] & b[15];
  wire p_15_0;
  wire g_15_0;
  wire p_15_1;
  wire g_15_1;
  wire p_15_2;
  wire g_15_2;
  wire p_15_3;
  wire g_15_3;
  wire p_15_4;
  wire g_15_4;
  wire p_15_5;
  wire g_15_5;
  wire p_15_6;
  wire g_15_6;
  wire p_15_7;
  wire g_15_7;
  wire p_15_8;
  wire g_15_8;
  wire p_15_9;
  wire g_15_9;
  wire p_15_10;
  wire g_15_10;
  wire p_15_11;
  wire g_15_11;
  wire p_15_12;
  wire g_15_12;
  wire p_15_13;
  wire g_15_13;
  wire p_15_14;
  wire g_15_14;
 assign sum[0] = p_0_0;
 assign p_1_0 = p_1_1 & p_0_0;
 assign g_1_0 = g_1_1 | (p_1_1 & g_0_0);
 assign sum[1] = p_1_1^ g_0_0;
 assign p_2_0 = p_2_1 & p_0_0;
 assign g_2_0 = g_2_1 | (p_2_1 & g_0_0);
 assign p_2_1 = p_2_2 & p_1_1;
 assign g_2_1 = g_2_2 | (p_2_2 & g_1_1);
 assign sum[2] = p_2_2^ g_1_0;
 assign p_3_0 = p_3_2 & p_1_0;
 assign g_3_0 = g_3_2 | (p_3_2 & g_1_0);
 assign p_3_1 = p_3_2 & p_1_1;
 assign g_3_1 = g_3_2 | (p_3_2 & g_1_1);
 assign p_3_2 = p_3_3 & p_2_2;
 assign g_3_2 = g_3_3 | (p_3_3 & g_2_2);
 assign sum[3] = p_3_3^ g_2_0;
 assign p_4_0 = p_4_1 & p_0_0;
 assign g_4_0 = g_4_1 | (p_4_1 & g_0_0);
 assign p_4_1 = p_4_3 & p_2_1;
 assign g_4_1 = g_4_3 | (p_4_3 & g_2_1);
 assign p_4_2 = p_4_3 & p_2_2;
 assign g_4_2 = g_4_3 | (p_4_3 & g_2_2);
 assign p_4_3 = p_4_4 & p_3_3;
 assign g_4_3 = g_4_4 | (p_4_4 & g_3_3);
 assign sum[4] = p_4_4^ g_3_0;
 assign p_5_0 = p_5_2 & p_1_0;
 assign g_5_0 = g_5_2 | (p_5_2 & g_1_0);
 assign p_5_1 = p_5_2 & p_1_1;
 assign g_5_1 = g_5_2 | (p_5_2 & g_1_1);
 assign p_5_2 = p_5_4 & p_3_2;
 assign g_5_2 = g_5_4 | (p_5_4 & g_3_2);
 assign p_5_3 = p_5_4 & p_3_3;
 assign g_5_3 = g_5_4 | (p_5_4 & g_3_3);
 assign p_5_4 = p_5_5 & p_4_4;
 assign g_5_4 = g_5_5 | (p_5_5 & g_4_4);
 assign sum[5] = p_5_5^ g_4_0;
 assign p_6_0 = p_6_3 & p_2_0;
 assign g_6_0 = g_6_3 | (p_6_3 & g_2_0);
 assign p_6_1 = p_6_3 & p_2_1;
 assign g_6_1 = g_6_3 | (p_6_3 & g_2_1);
 assign p_6_2 = p_6_3 & p_2_2;
 assign g_6_2 = g_6_3 | (p_6_3 & g_2_2);
 assign p_6_3 = p_6_5 & p_4_3;
 assign g_6_3 = g_6_5 | (p_6_5 & g_4_3);
 assign p_6_4 = p_6_5 & p_4_4;
 assign g_6_4 = g_6_5 | (p_6_5 & g_4_4);
 assign p_6_5 = p_6_6 & p_5_5;
 assign g_6_5 = g_6_6 | (p_6_6 & g_5_5);
 assign sum[6] = p_6_6^ g_5_0;
 assign p_7_0 = p_7_4 & p_3_0;
 assign g_7_0 = g_7_4 | (p_7_4 & g_3_0);
 assign p_7_1 = p_7_4 & p_3_1;
 assign g_7_1 = g_7_4 | (p_7_4 & g_3_1);
 assign p_7_2 = p_7_4 & p_3_2;
 assign g_7_2 = g_7_4 | (p_7_4 & g_3_2);
 assign p_7_3 = p_7_4 & p_3_3;
 assign g_7_3 = g_7_4 | (p_7_4 & g_3_3);
 assign p_7_4 = p_7_6 & p_5_4;
 assign g_7_4 = g_7_6 | (p_7_6 & g_5_4);
 assign p_7_5 = p_7_6 & p_5_5;
 assign g_7_5 = g_7_6 | (p_7_6 & g_5_5);
 assign p_7_6 = p_7_7 & p_6_6;
 assign g_7_6 = g_7_7 | (p_7_7 & g_6_6);
 assign sum[7] = p_7_7^ g_6_0;
 assign p_8_0 = p_8_1 & p_0_0;
 assign g_8_0 = g_8_1 | (p_8_1 & g_0_0);
 assign p_8_1 = p_8_5 & p_4_1;
 assign g_8_1 = g_8_5 | (p_8_5 & g_4_1);
 assign p_8_2 = p_8_5 & p_4_2;
 assign g_8_2 = g_8_5 | (p_8_5 & g_4_2);
 assign p_8_3 = p_8_5 & p_4_3;
 assign g_8_3 = g_8_5 | (p_8_5 & g_4_3);
 assign p_8_4 = p_8_5 & p_4_4;
 assign g_8_4 = g_8_5 | (p_8_5 & g_4_4);
 assign p_8_5 = p_8_7 & p_6_5;
 assign g_8_5 = g_8_7 | (p_8_7 & g_6_5);
 assign p_8_6 = p_8_7 & p_6_6;
 assign g_8_6 = g_8_7 | (p_8_7 & g_6_6);
 assign p_8_7 = p_8_8 & p_7_7;
 assign g_8_7 = g_8_8 | (p_8_8 & g_7_7);
 assign sum[8] = p_8_8^ g_7_0;
 assign p_9_0 = p_9_2 & p_1_0;
 assign g_9_0 = g_9_2 | (p_9_2 & g_1_0);
 assign p_9_1 = p_9_2 & p_1_1;
 assign g_9_1 = g_9_2 | (p_9_2 & g_1_1);
 assign p_9_2 = p_9_6 & p_5_2;
 assign g_9_2 = g_9_6 | (p_9_6 & g_5_2);
 assign p_9_3 = p_9_6 & p_5_3;
 assign g_9_3 = g_9_6 | (p_9_6 & g_5_3);
 assign p_9_4 = p_9_6 & p_5_4;
 assign g_9_4 = g_9_6 | (p_9_6 & g_5_4);
 assign p_9_5 = p_9_6 & p_5_5;
 assign g_9_5 = g_9_6 | (p_9_6 & g_5_5);
 assign p_9_6 = p_9_8 & p_7_6;
 assign g_9_6 = g_9_8 | (p_9_8 & g_7_6);
 assign p_9_7 = p_9_8 & p_7_7;
 assign g_9_7 = g_9_8 | (p_9_8 & g_7_7);
 assign p_9_8 = p_9_9 & p_8_8;
 assign g_9_8 = g_9_9 | (p_9_9 & g_8_8);
 assign sum[9] = p_9_9^ g_8_0;
 assign p_10_0 = p_10_3 & p_2_0;
 assign g_10_0 = g_10_3 | (p_10_3 & g_2_0);
 assign p_10_1 = p_10_3 & p_2_1;
 assign g_10_1 = g_10_3 | (p_10_3 & g_2_1);
 assign p_10_2 = p_10_3 & p_2_2;
 assign g_10_2 = g_10_3 | (p_10_3 & g_2_2);
 assign p_10_3 = p_10_7 & p_6_3;
 assign g_10_3 = g_10_7 | (p_10_7 & g_6_3);
 assign p_10_4 = p_10_7 & p_6_4;
 assign g_10_4 = g_10_7 | (p_10_7 & g_6_4);
 assign p_10_5 = p_10_7 & p_6_5;
 assign g_10_5 = g_10_7 | (p_10_7 & g_6_5);
 assign p_10_6 = p_10_7 & p_6_6;
 assign g_10_6 = g_10_7 | (p_10_7 & g_6_6);
 assign p_10_7 = p_10_9 & p_8_7;
 assign g_10_7 = g_10_9 | (p_10_9 & g_8_7);
 assign p_10_8 = p_10_9 & p_8_8;
 assign g_10_8 = g_10_9 | (p_10_9 & g_8_8);
 assign p_10_9 = p_10_10 & p_9_9;
 assign g_10_9 = g_10_10 | (p_10_10 & g_9_9);
 assign sum[10] = p_10_10^ g_9_0;
 assign p_11_0 = p_11_4 & p_3_0;
 assign g_11_0 = g_11_4 | (p_11_4 & g_3_0);
 assign p_11_1 = p_11_4 & p_3_1;
 assign g_11_1 = g_11_4 | (p_11_4 & g_3_1);
 assign p_11_2 = p_11_4 & p_3_2;
 assign g_11_2 = g_11_4 | (p_11_4 & g_3_2);
 assign p_11_3 = p_11_4 & p_3_3;
 assign g_11_3 = g_11_4 | (p_11_4 & g_3_3);
 assign p_11_4 = p_11_8 & p_7_4;
 assign g_11_4 = g_11_8 | (p_11_8 & g_7_4);
 assign p_11_5 = p_11_8 & p_7_5;
 assign g_11_5 = g_11_8 | (p_11_8 & g_7_5);
 assign p_11_6 = p_11_8 & p_7_6;
 assign g_11_6 = g_11_8 | (p_11_8 & g_7_6);
 assign p_11_7 = p_11_8 & p_7_7;
 assign g_11_7 = g_11_8 | (p_11_8 & g_7_7);
 assign p_11_8 = p_11_10 & p_9_8;
 assign g_11_8 = g_11_10 | (p_11_10 & g_9_8);
 assign p_11_9 = p_11_10 & p_9_9;
 assign g_11_9 = g_11_10 | (p_11_10 & g_9_9);
 assign p_11_10 = p_11_11 & p_10_10;
 assign g_11_10 = g_11_11 | (p_11_11 & g_10_10);
 assign sum[11] = p_11_11^ g_10_0;
 assign p_12_0 = p_12_5 & p_4_0;
 assign g_12_0 = g_12_5 | (p_12_5 & g_4_0);
 assign p_12_1 = p_12_5 & p_4_1;
 assign g_12_1 = g_12_5 | (p_12_5 & g_4_1);
 assign p_12_2 = p_12_5 & p_4_2;
 assign g_12_2 = g_12_5 | (p_12_5 & g_4_2);
 assign p_12_3 = p_12_5 & p_4_3;
 assign g_12_3 = g_12_5 | (p_12_5 & g_4_3);
 assign p_12_4 = p_12_5 & p_4_4;
 assign g_12_4 = g_12_5 | (p_12_5 & g_4_4);
 assign p_12_5 = p_12_9 & p_8_5;
 assign g_12_5 = g_12_9 | (p_12_9 & g_8_5);
 assign p_12_6 = p_12_9 & p_8_6;
 assign g_12_6 = g_12_9 | (p_12_9 & g_8_6);
 assign p_12_7 = p_12_9 & p_8_7;
 assign g_12_7 = g_12_9 | (p_12_9 & g_8_7);
 assign p_12_8 = p_12_9 & p_8_8;
 assign g_12_8 = g_12_9 | (p_12_9 & g_8_8);
 assign p_12_9 = p_12_11 & p_10_9;
 assign g_12_9 = g_12_11 | (p_12_11 & g_10_9);
 assign p_12_10 = p_12_11 & p_10_10;
 assign g_12_10 = g_12_11 | (p_12_11 & g_10_10);
 assign p_12_11 = p_12_12 & p_11_11;
 assign g_12_11 = g_12_12 | (p_12_12 & g_11_11);
 assign sum[12] = p_12_12^ g_11_0;
 assign p_13_0 = p_13_6 & p_5_0;
 assign g_13_0 = g_13_6 | (p_13_6 & g_5_0);
 assign p_13_1 = p_13_6 & p_5_1;
 assign g_13_1 = g_13_6 | (p_13_6 & g_5_1);
 assign p_13_2 = p_13_6 & p_5_2;
 assign g_13_2 = g_13_6 | (p_13_6 & g_5_2);
 assign p_13_3 = p_13_6 & p_5_3;
 assign g_13_3 = g_13_6 | (p_13_6 & g_5_3);
 assign p_13_4 = p_13_6 & p_5_4;
 assign g_13_4 = g_13_6 | (p_13_6 & g_5_4);
 assign p_13_5 = p_13_6 & p_5_5;
 assign g_13_5 = g_13_6 | (p_13_6 & g_5_5);
 assign p_13_6 = p_13_10 & p_9_6;
 assign g_13_6 = g_13_10 | (p_13_10 & g_9_6);
 assign p_13_7 = p_13_10 & p_9_7;
 assign g_13_7 = g_13_10 | (p_13_10 & g_9_7);
 assign p_13_8 = p_13_10 & p_9_8;
 assign g_13_8 = g_13_10 | (p_13_10 & g_9_8);
 assign p_13_9 = p_13_10 & p_9_9;
 assign g_13_9 = g_13_10 | (p_13_10 & g_9_9);
 assign p_13_10 = p_13_12 & p_11_10;
 assign g_13_10 = g_13_12 | (p_13_12 & g_11_10);
 assign p_13_11 = p_13_12 & p_11_11;
 assign g_13_11 = g_13_12 | (p_13_12 & g_11_11);
 assign p_13_12 = p_13_13 & p_12_12;
 assign g_13_12 = g_13_13 | (p_13_13 & g_12_12);
 assign sum[13] = p_13_13^ g_12_0;
 assign p_14_0 = p_14_7 & p_6_0;
 assign g_14_0 = g_14_7 | (p_14_7 & g_6_0);
 assign p_14_1 = p_14_7 & p_6_1;
 assign g_14_1 = g_14_7 | (p_14_7 & g_6_1);
 assign p_14_2 = p_14_7 & p_6_2;
 assign g_14_2 = g_14_7 | (p_14_7 & g_6_2);
 assign p_14_3 = p_14_7 & p_6_3;
 assign g_14_3 = g_14_7 | (p_14_7 & g_6_3);
 assign p_14_4 = p_14_7 & p_6_4;
 assign g_14_4 = g_14_7 | (p_14_7 & g_6_4);
 assign p_14_5 = p_14_7 & p_6_5;
 assign g_14_5 = g_14_7 | (p_14_7 & g_6_5);
 assign p_14_6 = p_14_7 & p_6_6;
 assign g_14_6 = g_14_7 | (p_14_7 & g_6_6);
 assign p_14_7 = p_14_11 & p_10_7;
 assign g_14_7 = g_14_11 | (p_14_11 & g_10_7);
 assign p_14_8 = p_14_11 & p_10_8;
 assign g_14_8 = g_14_11 | (p_14_11 & g_10_8);
 assign p_14_9 = p_14_11 & p_10_9;
 assign g_14_9 = g_14_11 | (p_14_11 & g_10_9);
 assign p_14_10 = p_14_11 & p_10_10;
 assign g_14_10 = g_14_11 | (p_14_11 & g_10_10);
 assign p_14_11 = p_14_13 & p_12_11;
 assign g_14_11 = g_14_13 | (p_14_13 & g_12_11);
 assign p_14_12 = p_14_13 & p_12_12;
 assign g_14_12 = g_14_13 | (p_14_13 & g_12_12);
 assign p_14_13 = p_14_14 & p_13_13;
 assign g_14_13 = g_14_14 | (p_14_14 & g_13_13);
 assign sum[14] = p_14_14^ g_13_0;
 assign p_15_0 = p_15_8 & p_7_0;
 assign g_15_0 = g_15_8 | (p_15_8 & g_7_0);
 assign p_15_1 = p_15_8 & p_7_1;
 assign g_15_1 = g_15_8 | (p_15_8 & g_7_1);
 assign p_15_2 = p_15_8 & p_7_2;
 assign g_15_2 = g_15_8 | (p_15_8 & g_7_2);
 assign p_15_3 = p_15_8 & p_7_3;
 assign g_15_3 = g_15_8 | (p_15_8 & g_7_3);
 assign p_15_4 = p_15_8 & p_7_4;
 assign g_15_4 = g_15_8 | (p_15_8 & g_7_4);
 assign p_15_5 = p_15_8 & p_7_5;
 assign g_15_5 = g_15_8 | (p_15_8 & g_7_5);
 assign p_15_6 = p_15_8 & p_7_6;
 assign g_15_6 = g_15_8 | (p_15_8 & g_7_6);
 assign p_15_7 = p_15_8 & p_7_7;
 assign g_15_7 = g_15_8 | (p_15_8 & g_7_7);
 assign p_15_8 = p_15_12 & p_11_8;
 assign g_15_8 = g_15_12 | (p_15_12 & g_11_8);
 assign p_15_9 = p_15_12 & p_11_9;
 assign g_15_9 = g_15_12 | (p_15_12 & g_11_9);
 assign p_15_10 = p_15_12 & p_11_10;
 assign g_15_10 = g_15_12 | (p_15_12 & g_11_10);
 assign p_15_11 = p_15_12 & p_11_11;
 assign g_15_11 = g_15_12 | (p_15_12 & g_11_11);
 assign p_15_12 = p_15_14 & p_13_12;
 assign g_15_12 = g_15_14 | (p_15_14 & g_13_12);
 assign p_15_13 = p_15_14 & p_13_13;
 assign g_15_13 = g_15_14 | (p_15_14 & g_13_13);
 assign p_15_14 = p_15_15 & p_14_14;
 assign g_15_14 = g_15_15 | (p_15_15 & g_14_14);
 assign sum[15] = p_15_15^ g_14_0;
 assign cout = g_15_0;
endmodule
