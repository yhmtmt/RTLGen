module MG_CPA(
  input [62:0] a,
  input [62:0] b,
  output [62:0] sum,
  output cout
);

  wire p_0_0;
  wire g_0_0;
 assign p_0_0 = a[0] ^ b[0];
 assign g_0_0 = a[0] & b[0];
  wire p_1_1;
  wire g_1_1;
 assign p_1_1 = a[1] ^ b[1];
 assign g_1_1 = a[1] & b[1];
  wire p_1_0;
  wire g_1_0;
  wire p_2_2;
  wire g_2_2;
 assign p_2_2 = a[2] ^ b[2];
 assign g_2_2 = a[2] & b[2];
  wire p_2_0;
  wire g_2_0;
  wire p_3_3;
  wire g_3_3;
 assign p_3_3 = a[3] ^ b[3];
 assign g_3_3 = a[3] & b[3];
  wire p_3_0;
  wire g_3_0;
  wire p_3_2;
  wire g_3_2;
  wire p_4_4;
  wire g_4_4;
 assign p_4_4 = a[4] ^ b[4];
 assign g_4_4 = a[4] & b[4];
  wire p_4_0;
  wire g_4_0;
  wire p_5_5;
  wire g_5_5;
 assign p_5_5 = a[5] ^ b[5];
 assign g_5_5 = a[5] & b[5];
  wire p_5_0;
  wire g_5_0;
  wire p_5_4;
  wire g_5_4;
  wire p_6_6;
  wire g_6_6;
 assign p_6_6 = a[6] ^ b[6];
 assign g_6_6 = a[6] & b[6];
  wire p_6_0;
  wire g_6_0;
  wire p_6_4;
  wire g_6_4;
  wire p_7_7;
  wire g_7_7;
 assign p_7_7 = a[7] ^ b[7];
 assign g_7_7 = a[7] & b[7];
  wire p_7_0;
  wire g_7_0;
  wire p_7_4;
  wire g_7_4;
  wire p_7_6;
  wire g_7_6;
  wire p_8_8;
  wire g_8_8;
 assign p_8_8 = a[8] ^ b[8];
 assign g_8_8 = a[8] & b[8];
  wire p_8_0;
  wire g_8_0;
  wire p_9_9;
  wire g_9_9;
 assign p_9_9 = a[9] ^ b[9];
 assign g_9_9 = a[9] & b[9];
  wire p_9_0;
  wire g_9_0;
  wire p_9_8;
  wire g_9_8;
  wire p_10_10;
  wire g_10_10;
 assign p_10_10 = a[10] ^ b[10];
 assign g_10_10 = a[10] & b[10];
  wire p_10_0;
  wire g_10_0;
  wire p_10_8;
  wire g_10_8;
  wire p_11_11;
  wire g_11_11;
 assign p_11_11 = a[11] ^ b[11];
 assign g_11_11 = a[11] & b[11];
  wire p_11_0;
  wire g_11_0;
  wire p_11_8;
  wire g_11_8;
  wire p_11_10;
  wire g_11_10;
  wire p_12_12;
  wire g_12_12;
 assign p_12_12 = a[12] ^ b[12];
 assign g_12_12 = a[12] & b[12];
  wire p_12_0;
  wire g_12_0;
  wire p_12_8;
  wire g_12_8;
  wire p_13_13;
  wire g_13_13;
 assign p_13_13 = a[13] ^ b[13];
 assign g_13_13 = a[13] & b[13];
  wire p_13_0;
  wire g_13_0;
  wire p_13_8;
  wire g_13_8;
  wire p_13_12;
  wire g_13_12;
  wire p_14_14;
  wire g_14_14;
 assign p_14_14 = a[14] ^ b[14];
 assign g_14_14 = a[14] & b[14];
  wire p_14_0;
  wire g_14_0;
  wire p_14_8;
  wire g_14_8;
  wire p_14_12;
  wire g_14_12;
  wire p_15_15;
  wire g_15_15;
 assign p_15_15 = a[15] ^ b[15];
 assign g_15_15 = a[15] & b[15];
  wire p_15_0;
  wire g_15_0;
  wire p_15_8;
  wire g_15_8;
  wire p_15_12;
  wire g_15_12;
  wire p_15_14;
  wire g_15_14;
  wire p_16_16;
  wire g_16_16;
 assign p_16_16 = a[16] ^ b[16];
 assign g_16_16 = a[16] & b[16];
  wire p_16_0;
  wire g_16_0;
  wire p_17_17;
  wire g_17_17;
 assign p_17_17 = a[17] ^ b[17];
 assign g_17_17 = a[17] & b[17];
  wire p_17_0;
  wire g_17_0;
  wire p_17_16;
  wire g_17_16;
  wire p_18_18;
  wire g_18_18;
 assign p_18_18 = a[18] ^ b[18];
 assign g_18_18 = a[18] & b[18];
  wire p_18_0;
  wire g_18_0;
  wire p_18_16;
  wire g_18_16;
  wire p_19_19;
  wire g_19_19;
 assign p_19_19 = a[19] ^ b[19];
 assign g_19_19 = a[19] & b[19];
  wire p_19_0;
  wire g_19_0;
  wire p_19_16;
  wire g_19_16;
  wire p_19_18;
  wire g_19_18;
  wire p_20_20;
  wire g_20_20;
 assign p_20_20 = a[20] ^ b[20];
 assign g_20_20 = a[20] & b[20];
  wire p_20_0;
  wire g_20_0;
  wire p_20_16;
  wire g_20_16;
  wire p_21_21;
  wire g_21_21;
 assign p_21_21 = a[21] ^ b[21];
 assign g_21_21 = a[21] & b[21];
  wire p_21_0;
  wire g_21_0;
  wire p_21_16;
  wire g_21_16;
  wire p_21_20;
  wire g_21_20;
  wire p_22_22;
  wire g_22_22;
 assign p_22_22 = a[22] ^ b[22];
 assign g_22_22 = a[22] & b[22];
  wire p_22_0;
  wire g_22_0;
  wire p_22_16;
  wire g_22_16;
  wire p_22_20;
  wire g_22_20;
  wire p_23_23;
  wire g_23_23;
 assign p_23_23 = a[23] ^ b[23];
 assign g_23_23 = a[23] & b[23];
  wire p_23_0;
  wire g_23_0;
  wire p_23_16;
  wire g_23_16;
  wire p_23_20;
  wire g_23_20;
  wire p_23_22;
  wire g_23_22;
  wire p_24_24;
  wire g_24_24;
 assign p_24_24 = a[24] ^ b[24];
 assign g_24_24 = a[24] & b[24];
  wire p_24_0;
  wire g_24_0;
  wire p_24_16;
  wire g_24_16;
  wire p_25_25;
  wire g_25_25;
 assign p_25_25 = a[25] ^ b[25];
 assign g_25_25 = a[25] & b[25];
  wire p_25_0;
  wire g_25_0;
  wire p_25_16;
  wire g_25_16;
  wire p_25_24;
  wire g_25_24;
  wire p_26_26;
  wire g_26_26;
 assign p_26_26 = a[26] ^ b[26];
 assign g_26_26 = a[26] & b[26];
  wire p_26_0;
  wire g_26_0;
  wire p_26_16;
  wire g_26_16;
  wire p_26_24;
  wire g_26_24;
  wire p_27_27;
  wire g_27_27;
 assign p_27_27 = a[27] ^ b[27];
 assign g_27_27 = a[27] & b[27];
  wire p_27_0;
  wire g_27_0;
  wire p_27_16;
  wire g_27_16;
  wire p_27_24;
  wire g_27_24;
  wire p_27_26;
  wire g_27_26;
  wire p_28_28;
  wire g_28_28;
 assign p_28_28 = a[28] ^ b[28];
 assign g_28_28 = a[28] & b[28];
  wire p_28_0;
  wire g_28_0;
  wire p_28_16;
  wire g_28_16;
  wire p_28_24;
  wire g_28_24;
  wire p_29_29;
  wire g_29_29;
 assign p_29_29 = a[29] ^ b[29];
 assign g_29_29 = a[29] & b[29];
  wire p_29_0;
  wire g_29_0;
  wire p_29_16;
  wire g_29_16;
  wire p_29_24;
  wire g_29_24;
  wire p_29_28;
  wire g_29_28;
  wire p_30_30;
  wire g_30_30;
 assign p_30_30 = a[30] ^ b[30];
 assign g_30_30 = a[30] & b[30];
  wire p_30_0;
  wire g_30_0;
  wire p_30_16;
  wire g_30_16;
  wire p_30_24;
  wire g_30_24;
  wire p_30_28;
  wire g_30_28;
  wire p_31_31;
  wire g_31_31;
 assign p_31_31 = a[31] ^ b[31];
 assign g_31_31 = a[31] & b[31];
  wire p_31_0;
  wire g_31_0;
  wire p_31_16;
  wire g_31_16;
  wire p_31_24;
  wire g_31_24;
  wire p_31_28;
  wire g_31_28;
  wire p_31_30;
  wire g_31_30;
  wire p_32_32;
  wire g_32_32;
 assign p_32_32 = a[32] ^ b[32];
 assign g_32_32 = a[32] & b[32];
  wire p_32_0;
  wire g_32_0;
  wire p_33_33;
  wire g_33_33;
 assign p_33_33 = a[33] ^ b[33];
 assign g_33_33 = a[33] & b[33];
  wire p_33_0;
  wire g_33_0;
  wire p_33_32;
  wire g_33_32;
  wire p_34_34;
  wire g_34_34;
 assign p_34_34 = a[34] ^ b[34];
 assign g_34_34 = a[34] & b[34];
  wire p_34_0;
  wire g_34_0;
  wire p_34_32;
  wire g_34_32;
  wire p_35_35;
  wire g_35_35;
 assign p_35_35 = a[35] ^ b[35];
 assign g_35_35 = a[35] & b[35];
  wire p_35_0;
  wire g_35_0;
  wire p_35_32;
  wire g_35_32;
  wire p_35_34;
  wire g_35_34;
  wire p_36_36;
  wire g_36_36;
 assign p_36_36 = a[36] ^ b[36];
 assign g_36_36 = a[36] & b[36];
  wire p_36_0;
  wire g_36_0;
  wire p_36_32;
  wire g_36_32;
  wire p_37_37;
  wire g_37_37;
 assign p_37_37 = a[37] ^ b[37];
 assign g_37_37 = a[37] & b[37];
  wire p_37_0;
  wire g_37_0;
  wire p_37_32;
  wire g_37_32;
  wire p_37_36;
  wire g_37_36;
  wire p_38_38;
  wire g_38_38;
 assign p_38_38 = a[38] ^ b[38];
 assign g_38_38 = a[38] & b[38];
  wire p_38_0;
  wire g_38_0;
  wire p_38_32;
  wire g_38_32;
  wire p_38_36;
  wire g_38_36;
  wire p_39_39;
  wire g_39_39;
 assign p_39_39 = a[39] ^ b[39];
 assign g_39_39 = a[39] & b[39];
  wire p_39_0;
  wire g_39_0;
  wire p_39_32;
  wire g_39_32;
  wire p_39_36;
  wire g_39_36;
  wire p_39_38;
  wire g_39_38;
  wire p_40_40;
  wire g_40_40;
 assign p_40_40 = a[40] ^ b[40];
 assign g_40_40 = a[40] & b[40];
  wire p_40_0;
  wire g_40_0;
  wire p_40_32;
  wire g_40_32;
  wire p_41_41;
  wire g_41_41;
 assign p_41_41 = a[41] ^ b[41];
 assign g_41_41 = a[41] & b[41];
  wire p_41_0;
  wire g_41_0;
  wire p_41_32;
  wire g_41_32;
  wire p_41_40;
  wire g_41_40;
  wire p_42_42;
  wire g_42_42;
 assign p_42_42 = a[42] ^ b[42];
 assign g_42_42 = a[42] & b[42];
  wire p_42_0;
  wire g_42_0;
  wire p_42_32;
  wire g_42_32;
  wire p_42_40;
  wire g_42_40;
  wire p_43_43;
  wire g_43_43;
 assign p_43_43 = a[43] ^ b[43];
 assign g_43_43 = a[43] & b[43];
  wire p_43_0;
  wire g_43_0;
  wire p_43_32;
  wire g_43_32;
  wire p_43_40;
  wire g_43_40;
  wire p_43_42;
  wire g_43_42;
  wire p_44_44;
  wire g_44_44;
 assign p_44_44 = a[44] ^ b[44];
 assign g_44_44 = a[44] & b[44];
  wire p_44_0;
  wire g_44_0;
  wire p_44_32;
  wire g_44_32;
  wire p_44_40;
  wire g_44_40;
  wire p_45_45;
  wire g_45_45;
 assign p_45_45 = a[45] ^ b[45];
 assign g_45_45 = a[45] & b[45];
  wire p_45_0;
  wire g_45_0;
  wire p_45_32;
  wire g_45_32;
  wire p_45_40;
  wire g_45_40;
  wire p_45_44;
  wire g_45_44;
  wire p_46_46;
  wire g_46_46;
 assign p_46_46 = a[46] ^ b[46];
 assign g_46_46 = a[46] & b[46];
  wire p_46_0;
  wire g_46_0;
  wire p_46_32;
  wire g_46_32;
  wire p_46_40;
  wire g_46_40;
  wire p_46_44;
  wire g_46_44;
  wire p_47_47;
  wire g_47_47;
 assign p_47_47 = a[47] ^ b[47];
 assign g_47_47 = a[47] & b[47];
  wire p_47_0;
  wire g_47_0;
  wire p_47_32;
  wire g_47_32;
  wire p_47_40;
  wire g_47_40;
  wire p_47_44;
  wire g_47_44;
  wire p_47_46;
  wire g_47_46;
  wire p_48_48;
  wire g_48_48;
 assign p_48_48 = a[48] ^ b[48];
 assign g_48_48 = a[48] & b[48];
  wire p_48_0;
  wire g_48_0;
  wire p_48_32;
  wire g_48_32;
  wire p_49_49;
  wire g_49_49;
 assign p_49_49 = a[49] ^ b[49];
 assign g_49_49 = a[49] & b[49];
  wire p_49_0;
  wire g_49_0;
  wire p_49_32;
  wire g_49_32;
  wire p_49_48;
  wire g_49_48;
  wire p_50_50;
  wire g_50_50;
 assign p_50_50 = a[50] ^ b[50];
 assign g_50_50 = a[50] & b[50];
  wire p_50_0;
  wire g_50_0;
  wire p_50_32;
  wire g_50_32;
  wire p_50_48;
  wire g_50_48;
  wire p_51_51;
  wire g_51_51;
 assign p_51_51 = a[51] ^ b[51];
 assign g_51_51 = a[51] & b[51];
  wire p_51_0;
  wire g_51_0;
  wire p_51_32;
  wire g_51_32;
  wire p_51_48;
  wire g_51_48;
  wire p_51_50;
  wire g_51_50;
  wire p_52_52;
  wire g_52_52;
 assign p_52_52 = a[52] ^ b[52];
 assign g_52_52 = a[52] & b[52];
  wire p_52_0;
  wire g_52_0;
  wire p_52_32;
  wire g_52_32;
  wire p_52_48;
  wire g_52_48;
  wire p_53_53;
  wire g_53_53;
 assign p_53_53 = a[53] ^ b[53];
 assign g_53_53 = a[53] & b[53];
  wire p_53_0;
  wire g_53_0;
  wire p_53_32;
  wire g_53_32;
  wire p_53_48;
  wire g_53_48;
  wire p_53_52;
  wire g_53_52;
  wire p_54_54;
  wire g_54_54;
 assign p_54_54 = a[54] ^ b[54];
 assign g_54_54 = a[54] & b[54];
  wire p_54_0;
  wire g_54_0;
  wire p_54_32;
  wire g_54_32;
  wire p_54_48;
  wire g_54_48;
  wire p_54_52;
  wire g_54_52;
  wire p_55_55;
  wire g_55_55;
 assign p_55_55 = a[55] ^ b[55];
 assign g_55_55 = a[55] & b[55];
  wire p_55_0;
  wire g_55_0;
  wire p_55_32;
  wire g_55_32;
  wire p_55_48;
  wire g_55_48;
  wire p_55_52;
  wire g_55_52;
  wire p_55_54;
  wire g_55_54;
  wire p_56_56;
  wire g_56_56;
 assign p_56_56 = a[56] ^ b[56];
 assign g_56_56 = a[56] & b[56];
  wire p_56_0;
  wire g_56_0;
  wire p_56_32;
  wire g_56_32;
  wire p_56_48;
  wire g_56_48;
  wire p_57_57;
  wire g_57_57;
 assign p_57_57 = a[57] ^ b[57];
 assign g_57_57 = a[57] & b[57];
  wire p_57_0;
  wire g_57_0;
  wire p_57_32;
  wire g_57_32;
  wire p_57_48;
  wire g_57_48;
  wire p_57_56;
  wire g_57_56;
  wire p_58_58;
  wire g_58_58;
 assign p_58_58 = a[58] ^ b[58];
 assign g_58_58 = a[58] & b[58];
  wire p_58_0;
  wire g_58_0;
  wire p_58_32;
  wire g_58_32;
  wire p_58_48;
  wire g_58_48;
  wire p_58_56;
  wire g_58_56;
  wire p_59_59;
  wire g_59_59;
 assign p_59_59 = a[59] ^ b[59];
 assign g_59_59 = a[59] & b[59];
  wire p_59_0;
  wire g_59_0;
  wire p_59_32;
  wire g_59_32;
  wire p_59_48;
  wire g_59_48;
  wire p_59_56;
  wire g_59_56;
  wire p_59_58;
  wire g_59_58;
  wire p_60_60;
  wire g_60_60;
 assign p_60_60 = a[60] ^ b[60];
 assign g_60_60 = a[60] & b[60];
  wire p_60_0;
  wire g_60_0;
  wire p_60_32;
  wire g_60_32;
  wire p_60_48;
  wire g_60_48;
  wire p_60_56;
  wire g_60_56;
  wire p_61_61;
  wire g_61_61;
 assign p_61_61 = a[61] ^ b[61];
 assign g_61_61 = a[61] & b[61];
  wire p_61_0;
  wire g_61_0;
  wire p_61_32;
  wire g_61_32;
  wire p_61_48;
  wire g_61_48;
  wire p_61_56;
  wire g_61_56;
  wire p_61_60;
  wire g_61_60;
  wire p_62_62;
  wire g_62_62;
 assign p_62_62 = a[62] ^ b[62];
 assign g_62_62 = a[62] & b[62];
  wire p_62_0;
  wire g_62_0;
  wire p_62_32;
  wire g_62_32;
  wire p_62_48;
  wire g_62_48;
  wire p_62_56;
  wire g_62_56;
  wire p_62_60;
  wire g_62_60;
 assign sum[0] = p_0_0;
 assign p_1_0 = p_1_1 & p_0_0;
 assign g_1_0 = g_1_1 | (p_1_1 & g_0_0);
 assign sum[1] = p_1_1^ g_0_0;
 assign p_2_0 = p_2_2 & p_1_0;
 assign g_2_0 = g_2_2 | (p_2_2 & g_1_0);
 assign sum[2] = p_2_2^ g_1_0;
 assign p_3_0 = p_3_2 & p_1_0;
 assign g_3_0 = g_3_2 | (p_3_2 & g_1_0);
 assign p_3_2 = p_3_3 & p_2_2;
 assign g_3_2 = g_3_3 | (p_3_3 & g_2_2);
 assign sum[3] = p_3_3^ g_2_0;
 assign p_4_0 = p_4_4 & p_3_0;
 assign g_4_0 = g_4_4 | (p_4_4 & g_3_0);
 assign sum[4] = p_4_4^ g_3_0;
 assign p_5_0 = p_5_4 & p_3_0;
 assign g_5_0 = g_5_4 | (p_5_4 & g_3_0);
 assign p_5_4 = p_5_5 & p_4_4;
 assign g_5_4 = g_5_5 | (p_5_5 & g_4_4);
 assign sum[5] = p_5_5^ g_4_0;
 assign p_6_0 = p_6_4 & p_3_0;
 assign g_6_0 = g_6_4 | (p_6_4 & g_3_0);
 assign p_6_4 = p_6_6 & p_5_4;
 assign g_6_4 = g_6_6 | (p_6_6 & g_5_4);
 assign sum[6] = p_6_6^ g_5_0;
 assign p_7_0 = p_7_4 & p_3_0;
 assign g_7_0 = g_7_4 | (p_7_4 & g_3_0);
 assign p_7_4 = p_7_6 & p_5_4;
 assign g_7_4 = g_7_6 | (p_7_6 & g_5_4);
 assign p_7_6 = p_7_7 & p_6_6;
 assign g_7_6 = g_7_7 | (p_7_7 & g_6_6);
 assign sum[7] = p_7_7^ g_6_0;
 assign p_8_0 = p_8_8 & p_7_0;
 assign g_8_0 = g_8_8 | (p_8_8 & g_7_0);
 assign sum[8] = p_8_8^ g_7_0;
 assign p_9_0 = p_9_8 & p_7_0;
 assign g_9_0 = g_9_8 | (p_9_8 & g_7_0);
 assign p_9_8 = p_9_9 & p_8_8;
 assign g_9_8 = g_9_9 | (p_9_9 & g_8_8);
 assign sum[9] = p_9_9^ g_8_0;
 assign p_10_0 = p_10_8 & p_7_0;
 assign g_10_0 = g_10_8 | (p_10_8 & g_7_0);
 assign p_10_8 = p_10_10 & p_9_8;
 assign g_10_8 = g_10_10 | (p_10_10 & g_9_8);
 assign sum[10] = p_10_10^ g_9_0;
 assign p_11_0 = p_11_8 & p_7_0;
 assign g_11_0 = g_11_8 | (p_11_8 & g_7_0);
 assign p_11_8 = p_11_10 & p_9_8;
 assign g_11_8 = g_11_10 | (p_11_10 & g_9_8);
 assign p_11_10 = p_11_11 & p_10_10;
 assign g_11_10 = g_11_11 | (p_11_11 & g_10_10);
 assign sum[11] = p_11_11^ g_10_0;
 assign p_12_0 = p_12_8 & p_7_0;
 assign g_12_0 = g_12_8 | (p_12_8 & g_7_0);
 assign p_12_8 = p_12_12 & p_11_8;
 assign g_12_8 = g_12_12 | (p_12_12 & g_11_8);
 assign sum[12] = p_12_12^ g_11_0;
 assign p_13_0 = p_13_8 & p_7_0;
 assign g_13_0 = g_13_8 | (p_13_8 & g_7_0);
 assign p_13_8 = p_13_12 & p_11_8;
 assign g_13_8 = g_13_12 | (p_13_12 & g_11_8);
 assign p_13_12 = p_13_13 & p_12_12;
 assign g_13_12 = g_13_13 | (p_13_13 & g_12_12);
 assign sum[13] = p_13_13^ g_12_0;
 assign p_14_0 = p_14_8 & p_7_0;
 assign g_14_0 = g_14_8 | (p_14_8 & g_7_0);
 assign p_14_8 = p_14_12 & p_11_8;
 assign g_14_8 = g_14_12 | (p_14_12 & g_11_8);
 assign p_14_12 = p_14_14 & p_13_12;
 assign g_14_12 = g_14_14 | (p_14_14 & g_13_12);
 assign sum[14] = p_14_14^ g_13_0;
 assign p_15_0 = p_15_8 & p_7_0;
 assign g_15_0 = g_15_8 | (p_15_8 & g_7_0);
 assign p_15_8 = p_15_12 & p_11_8;
 assign g_15_8 = g_15_12 | (p_15_12 & g_11_8);
 assign p_15_12 = p_15_14 & p_13_12;
 assign g_15_12 = g_15_14 | (p_15_14 & g_13_12);
 assign p_15_14 = p_15_15 & p_14_14;
 assign g_15_14 = g_15_15 | (p_15_15 & g_14_14);
 assign sum[15] = p_15_15^ g_14_0;
 assign p_16_0 = p_16_16 & p_15_0;
 assign g_16_0 = g_16_16 | (p_16_16 & g_15_0);
 assign sum[16] = p_16_16^ g_15_0;
 assign p_17_0 = p_17_16 & p_15_0;
 assign g_17_0 = g_17_16 | (p_17_16 & g_15_0);
 assign p_17_16 = p_17_17 & p_16_16;
 assign g_17_16 = g_17_17 | (p_17_17 & g_16_16);
 assign sum[17] = p_17_17^ g_16_0;
 assign p_18_0 = p_18_16 & p_15_0;
 assign g_18_0 = g_18_16 | (p_18_16 & g_15_0);
 assign p_18_16 = p_18_18 & p_17_16;
 assign g_18_16 = g_18_18 | (p_18_18 & g_17_16);
 assign sum[18] = p_18_18^ g_17_0;
 assign p_19_0 = p_19_16 & p_15_0;
 assign g_19_0 = g_19_16 | (p_19_16 & g_15_0);
 assign p_19_16 = p_19_18 & p_17_16;
 assign g_19_16 = g_19_18 | (p_19_18 & g_17_16);
 assign p_19_18 = p_19_19 & p_18_18;
 assign g_19_18 = g_19_19 | (p_19_19 & g_18_18);
 assign sum[19] = p_19_19^ g_18_0;
 assign p_20_0 = p_20_16 & p_15_0;
 assign g_20_0 = g_20_16 | (p_20_16 & g_15_0);
 assign p_20_16 = p_20_20 & p_19_16;
 assign g_20_16 = g_20_20 | (p_20_20 & g_19_16);
 assign sum[20] = p_20_20^ g_19_0;
 assign p_21_0 = p_21_16 & p_15_0;
 assign g_21_0 = g_21_16 | (p_21_16 & g_15_0);
 assign p_21_16 = p_21_20 & p_19_16;
 assign g_21_16 = g_21_20 | (p_21_20 & g_19_16);
 assign p_21_20 = p_21_21 & p_20_20;
 assign g_21_20 = g_21_21 | (p_21_21 & g_20_20);
 assign sum[21] = p_21_21^ g_20_0;
 assign p_22_0 = p_22_16 & p_15_0;
 assign g_22_0 = g_22_16 | (p_22_16 & g_15_0);
 assign p_22_16 = p_22_20 & p_19_16;
 assign g_22_16 = g_22_20 | (p_22_20 & g_19_16);
 assign p_22_20 = p_22_22 & p_21_20;
 assign g_22_20 = g_22_22 | (p_22_22 & g_21_20);
 assign sum[22] = p_22_22^ g_21_0;
 assign p_23_0 = p_23_16 & p_15_0;
 assign g_23_0 = g_23_16 | (p_23_16 & g_15_0);
 assign p_23_16 = p_23_20 & p_19_16;
 assign g_23_16 = g_23_20 | (p_23_20 & g_19_16);
 assign p_23_20 = p_23_22 & p_21_20;
 assign g_23_20 = g_23_22 | (p_23_22 & g_21_20);
 assign p_23_22 = p_23_23 & p_22_22;
 assign g_23_22 = g_23_23 | (p_23_23 & g_22_22);
 assign sum[23] = p_23_23^ g_22_0;
 assign p_24_0 = p_24_16 & p_15_0;
 assign g_24_0 = g_24_16 | (p_24_16 & g_15_0);
 assign p_24_16 = p_24_24 & p_23_16;
 assign g_24_16 = g_24_24 | (p_24_24 & g_23_16);
 assign sum[24] = p_24_24^ g_23_0;
 assign p_25_0 = p_25_16 & p_15_0;
 assign g_25_0 = g_25_16 | (p_25_16 & g_15_0);
 assign p_25_16 = p_25_24 & p_23_16;
 assign g_25_16 = g_25_24 | (p_25_24 & g_23_16);
 assign p_25_24 = p_25_25 & p_24_24;
 assign g_25_24 = g_25_25 | (p_25_25 & g_24_24);
 assign sum[25] = p_25_25^ g_24_0;
 assign p_26_0 = p_26_16 & p_15_0;
 assign g_26_0 = g_26_16 | (p_26_16 & g_15_0);
 assign p_26_16 = p_26_24 & p_23_16;
 assign g_26_16 = g_26_24 | (p_26_24 & g_23_16);
 assign p_26_24 = p_26_26 & p_25_24;
 assign g_26_24 = g_26_26 | (p_26_26 & g_25_24);
 assign sum[26] = p_26_26^ g_25_0;
 assign p_27_0 = p_27_16 & p_15_0;
 assign g_27_0 = g_27_16 | (p_27_16 & g_15_0);
 assign p_27_16 = p_27_24 & p_23_16;
 assign g_27_16 = g_27_24 | (p_27_24 & g_23_16);
 assign p_27_24 = p_27_26 & p_25_24;
 assign g_27_24 = g_27_26 | (p_27_26 & g_25_24);
 assign p_27_26 = p_27_27 & p_26_26;
 assign g_27_26 = g_27_27 | (p_27_27 & g_26_26);
 assign sum[27] = p_27_27^ g_26_0;
 assign p_28_0 = p_28_16 & p_15_0;
 assign g_28_0 = g_28_16 | (p_28_16 & g_15_0);
 assign p_28_16 = p_28_24 & p_23_16;
 assign g_28_16 = g_28_24 | (p_28_24 & g_23_16);
 assign p_28_24 = p_28_28 & p_27_24;
 assign g_28_24 = g_28_28 | (p_28_28 & g_27_24);
 assign sum[28] = p_28_28^ g_27_0;
 assign p_29_0 = p_29_16 & p_15_0;
 assign g_29_0 = g_29_16 | (p_29_16 & g_15_0);
 assign p_29_16 = p_29_24 & p_23_16;
 assign g_29_16 = g_29_24 | (p_29_24 & g_23_16);
 assign p_29_24 = p_29_28 & p_27_24;
 assign g_29_24 = g_29_28 | (p_29_28 & g_27_24);
 assign p_29_28 = p_29_29 & p_28_28;
 assign g_29_28 = g_29_29 | (p_29_29 & g_28_28);
 assign sum[29] = p_29_29^ g_28_0;
 assign p_30_0 = p_30_16 & p_15_0;
 assign g_30_0 = g_30_16 | (p_30_16 & g_15_0);
 assign p_30_16 = p_30_24 & p_23_16;
 assign g_30_16 = g_30_24 | (p_30_24 & g_23_16);
 assign p_30_24 = p_30_28 & p_27_24;
 assign g_30_24 = g_30_28 | (p_30_28 & g_27_24);
 assign p_30_28 = p_30_30 & p_29_28;
 assign g_30_28 = g_30_30 | (p_30_30 & g_29_28);
 assign sum[30] = p_30_30^ g_29_0;
 assign p_31_0 = p_31_16 & p_15_0;
 assign g_31_0 = g_31_16 | (p_31_16 & g_15_0);
 assign p_31_16 = p_31_24 & p_23_16;
 assign g_31_16 = g_31_24 | (p_31_24 & g_23_16);
 assign p_31_24 = p_31_28 & p_27_24;
 assign g_31_24 = g_31_28 | (p_31_28 & g_27_24);
 assign p_31_28 = p_31_30 & p_29_28;
 assign g_31_28 = g_31_30 | (p_31_30 & g_29_28);
 assign p_31_30 = p_31_31 & p_30_30;
 assign g_31_30 = g_31_31 | (p_31_31 & g_30_30);
 assign sum[31] = p_31_31^ g_30_0;
 assign p_32_0 = p_32_32 & p_31_0;
 assign g_32_0 = g_32_32 | (p_32_32 & g_31_0);
 assign sum[32] = p_32_32^ g_31_0;
 assign p_33_0 = p_33_32 & p_31_0;
 assign g_33_0 = g_33_32 | (p_33_32 & g_31_0);
 assign p_33_32 = p_33_33 & p_32_32;
 assign g_33_32 = g_33_33 | (p_33_33 & g_32_32);
 assign sum[33] = p_33_33^ g_32_0;
 assign p_34_0 = p_34_32 & p_31_0;
 assign g_34_0 = g_34_32 | (p_34_32 & g_31_0);
 assign p_34_32 = p_34_34 & p_33_32;
 assign g_34_32 = g_34_34 | (p_34_34 & g_33_32);
 assign sum[34] = p_34_34^ g_33_0;
 assign p_35_0 = p_35_32 & p_31_0;
 assign g_35_0 = g_35_32 | (p_35_32 & g_31_0);
 assign p_35_32 = p_35_34 & p_33_32;
 assign g_35_32 = g_35_34 | (p_35_34 & g_33_32);
 assign p_35_34 = p_35_35 & p_34_34;
 assign g_35_34 = g_35_35 | (p_35_35 & g_34_34);
 assign sum[35] = p_35_35^ g_34_0;
 assign p_36_0 = p_36_32 & p_31_0;
 assign g_36_0 = g_36_32 | (p_36_32 & g_31_0);
 assign p_36_32 = p_36_36 & p_35_32;
 assign g_36_32 = g_36_36 | (p_36_36 & g_35_32);
 assign sum[36] = p_36_36^ g_35_0;
 assign p_37_0 = p_37_32 & p_31_0;
 assign g_37_0 = g_37_32 | (p_37_32 & g_31_0);
 assign p_37_32 = p_37_36 & p_35_32;
 assign g_37_32 = g_37_36 | (p_37_36 & g_35_32);
 assign p_37_36 = p_37_37 & p_36_36;
 assign g_37_36 = g_37_37 | (p_37_37 & g_36_36);
 assign sum[37] = p_37_37^ g_36_0;
 assign p_38_0 = p_38_32 & p_31_0;
 assign g_38_0 = g_38_32 | (p_38_32 & g_31_0);
 assign p_38_32 = p_38_36 & p_35_32;
 assign g_38_32 = g_38_36 | (p_38_36 & g_35_32);
 assign p_38_36 = p_38_38 & p_37_36;
 assign g_38_36 = g_38_38 | (p_38_38 & g_37_36);
 assign sum[38] = p_38_38^ g_37_0;
 assign p_39_0 = p_39_32 & p_31_0;
 assign g_39_0 = g_39_32 | (p_39_32 & g_31_0);
 assign p_39_32 = p_39_36 & p_35_32;
 assign g_39_32 = g_39_36 | (p_39_36 & g_35_32);
 assign p_39_36 = p_39_38 & p_37_36;
 assign g_39_36 = g_39_38 | (p_39_38 & g_37_36);
 assign p_39_38 = p_39_39 & p_38_38;
 assign g_39_38 = g_39_39 | (p_39_39 & g_38_38);
 assign sum[39] = p_39_39^ g_38_0;
 assign p_40_0 = p_40_32 & p_31_0;
 assign g_40_0 = g_40_32 | (p_40_32 & g_31_0);
 assign p_40_32 = p_40_40 & p_39_32;
 assign g_40_32 = g_40_40 | (p_40_40 & g_39_32);
 assign sum[40] = p_40_40^ g_39_0;
 assign p_41_0 = p_41_32 & p_31_0;
 assign g_41_0 = g_41_32 | (p_41_32 & g_31_0);
 assign p_41_32 = p_41_40 & p_39_32;
 assign g_41_32 = g_41_40 | (p_41_40 & g_39_32);
 assign p_41_40 = p_41_41 & p_40_40;
 assign g_41_40 = g_41_41 | (p_41_41 & g_40_40);
 assign sum[41] = p_41_41^ g_40_0;
 assign p_42_0 = p_42_32 & p_31_0;
 assign g_42_0 = g_42_32 | (p_42_32 & g_31_0);
 assign p_42_32 = p_42_40 & p_39_32;
 assign g_42_32 = g_42_40 | (p_42_40 & g_39_32);
 assign p_42_40 = p_42_42 & p_41_40;
 assign g_42_40 = g_42_42 | (p_42_42 & g_41_40);
 assign sum[42] = p_42_42^ g_41_0;
 assign p_43_0 = p_43_32 & p_31_0;
 assign g_43_0 = g_43_32 | (p_43_32 & g_31_0);
 assign p_43_32 = p_43_40 & p_39_32;
 assign g_43_32 = g_43_40 | (p_43_40 & g_39_32);
 assign p_43_40 = p_43_42 & p_41_40;
 assign g_43_40 = g_43_42 | (p_43_42 & g_41_40);
 assign p_43_42 = p_43_43 & p_42_42;
 assign g_43_42 = g_43_43 | (p_43_43 & g_42_42);
 assign sum[43] = p_43_43^ g_42_0;
 assign p_44_0 = p_44_32 & p_31_0;
 assign g_44_0 = g_44_32 | (p_44_32 & g_31_0);
 assign p_44_32 = p_44_40 & p_39_32;
 assign g_44_32 = g_44_40 | (p_44_40 & g_39_32);
 assign p_44_40 = p_44_44 & p_43_40;
 assign g_44_40 = g_44_44 | (p_44_44 & g_43_40);
 assign sum[44] = p_44_44^ g_43_0;
 assign p_45_0 = p_45_32 & p_31_0;
 assign g_45_0 = g_45_32 | (p_45_32 & g_31_0);
 assign p_45_32 = p_45_40 & p_39_32;
 assign g_45_32 = g_45_40 | (p_45_40 & g_39_32);
 assign p_45_40 = p_45_44 & p_43_40;
 assign g_45_40 = g_45_44 | (p_45_44 & g_43_40);
 assign p_45_44 = p_45_45 & p_44_44;
 assign g_45_44 = g_45_45 | (p_45_45 & g_44_44);
 assign sum[45] = p_45_45^ g_44_0;
 assign p_46_0 = p_46_32 & p_31_0;
 assign g_46_0 = g_46_32 | (p_46_32 & g_31_0);
 assign p_46_32 = p_46_40 & p_39_32;
 assign g_46_32 = g_46_40 | (p_46_40 & g_39_32);
 assign p_46_40 = p_46_44 & p_43_40;
 assign g_46_40 = g_46_44 | (p_46_44 & g_43_40);
 assign p_46_44 = p_46_46 & p_45_44;
 assign g_46_44 = g_46_46 | (p_46_46 & g_45_44);
 assign sum[46] = p_46_46^ g_45_0;
 assign p_47_0 = p_47_32 & p_31_0;
 assign g_47_0 = g_47_32 | (p_47_32 & g_31_0);
 assign p_47_32 = p_47_40 & p_39_32;
 assign g_47_32 = g_47_40 | (p_47_40 & g_39_32);
 assign p_47_40 = p_47_44 & p_43_40;
 assign g_47_40 = g_47_44 | (p_47_44 & g_43_40);
 assign p_47_44 = p_47_46 & p_45_44;
 assign g_47_44 = g_47_46 | (p_47_46 & g_45_44);
 assign p_47_46 = p_47_47 & p_46_46;
 assign g_47_46 = g_47_47 | (p_47_47 & g_46_46);
 assign sum[47] = p_47_47^ g_46_0;
 assign p_48_0 = p_48_32 & p_31_0;
 assign g_48_0 = g_48_32 | (p_48_32 & g_31_0);
 assign p_48_32 = p_48_48 & p_47_32;
 assign g_48_32 = g_48_48 | (p_48_48 & g_47_32);
 assign sum[48] = p_48_48^ g_47_0;
 assign p_49_0 = p_49_32 & p_31_0;
 assign g_49_0 = g_49_32 | (p_49_32 & g_31_0);
 assign p_49_32 = p_49_48 & p_47_32;
 assign g_49_32 = g_49_48 | (p_49_48 & g_47_32);
 assign p_49_48 = p_49_49 & p_48_48;
 assign g_49_48 = g_49_49 | (p_49_49 & g_48_48);
 assign sum[49] = p_49_49^ g_48_0;
 assign p_50_0 = p_50_32 & p_31_0;
 assign g_50_0 = g_50_32 | (p_50_32 & g_31_0);
 assign p_50_32 = p_50_48 & p_47_32;
 assign g_50_32 = g_50_48 | (p_50_48 & g_47_32);
 assign p_50_48 = p_50_50 & p_49_48;
 assign g_50_48 = g_50_50 | (p_50_50 & g_49_48);
 assign sum[50] = p_50_50^ g_49_0;
 assign p_51_0 = p_51_32 & p_31_0;
 assign g_51_0 = g_51_32 | (p_51_32 & g_31_0);
 assign p_51_32 = p_51_48 & p_47_32;
 assign g_51_32 = g_51_48 | (p_51_48 & g_47_32);
 assign p_51_48 = p_51_50 & p_49_48;
 assign g_51_48 = g_51_50 | (p_51_50 & g_49_48);
 assign p_51_50 = p_51_51 & p_50_50;
 assign g_51_50 = g_51_51 | (p_51_51 & g_50_50);
 assign sum[51] = p_51_51^ g_50_0;
 assign p_52_0 = p_52_32 & p_31_0;
 assign g_52_0 = g_52_32 | (p_52_32 & g_31_0);
 assign p_52_32 = p_52_48 & p_47_32;
 assign g_52_32 = g_52_48 | (p_52_48 & g_47_32);
 assign p_52_48 = p_52_52 & p_51_48;
 assign g_52_48 = g_52_52 | (p_52_52 & g_51_48);
 assign sum[52] = p_52_52^ g_51_0;
 assign p_53_0 = p_53_32 & p_31_0;
 assign g_53_0 = g_53_32 | (p_53_32 & g_31_0);
 assign p_53_32 = p_53_48 & p_47_32;
 assign g_53_32 = g_53_48 | (p_53_48 & g_47_32);
 assign p_53_48 = p_53_52 & p_51_48;
 assign g_53_48 = g_53_52 | (p_53_52 & g_51_48);
 assign p_53_52 = p_53_53 & p_52_52;
 assign g_53_52 = g_53_53 | (p_53_53 & g_52_52);
 assign sum[53] = p_53_53^ g_52_0;
 assign p_54_0 = p_54_32 & p_31_0;
 assign g_54_0 = g_54_32 | (p_54_32 & g_31_0);
 assign p_54_32 = p_54_48 & p_47_32;
 assign g_54_32 = g_54_48 | (p_54_48 & g_47_32);
 assign p_54_48 = p_54_52 & p_51_48;
 assign g_54_48 = g_54_52 | (p_54_52 & g_51_48);
 assign p_54_52 = p_54_54 & p_53_52;
 assign g_54_52 = g_54_54 | (p_54_54 & g_53_52);
 assign sum[54] = p_54_54^ g_53_0;
 assign p_55_0 = p_55_32 & p_31_0;
 assign g_55_0 = g_55_32 | (p_55_32 & g_31_0);
 assign p_55_32 = p_55_48 & p_47_32;
 assign g_55_32 = g_55_48 | (p_55_48 & g_47_32);
 assign p_55_48 = p_55_52 & p_51_48;
 assign g_55_48 = g_55_52 | (p_55_52 & g_51_48);
 assign p_55_52 = p_55_54 & p_53_52;
 assign g_55_52 = g_55_54 | (p_55_54 & g_53_52);
 assign p_55_54 = p_55_55 & p_54_54;
 assign g_55_54 = g_55_55 | (p_55_55 & g_54_54);
 assign sum[55] = p_55_55^ g_54_0;
 assign p_56_0 = p_56_32 & p_31_0;
 assign g_56_0 = g_56_32 | (p_56_32 & g_31_0);
 assign p_56_32 = p_56_48 & p_47_32;
 assign g_56_32 = g_56_48 | (p_56_48 & g_47_32);
 assign p_56_48 = p_56_56 & p_55_48;
 assign g_56_48 = g_56_56 | (p_56_56 & g_55_48);
 assign sum[56] = p_56_56^ g_55_0;
 assign p_57_0 = p_57_32 & p_31_0;
 assign g_57_0 = g_57_32 | (p_57_32 & g_31_0);
 assign p_57_32 = p_57_48 & p_47_32;
 assign g_57_32 = g_57_48 | (p_57_48 & g_47_32);
 assign p_57_48 = p_57_56 & p_55_48;
 assign g_57_48 = g_57_56 | (p_57_56 & g_55_48);
 assign p_57_56 = p_57_57 & p_56_56;
 assign g_57_56 = g_57_57 | (p_57_57 & g_56_56);
 assign sum[57] = p_57_57^ g_56_0;
 assign p_58_0 = p_58_32 & p_31_0;
 assign g_58_0 = g_58_32 | (p_58_32 & g_31_0);
 assign p_58_32 = p_58_48 & p_47_32;
 assign g_58_32 = g_58_48 | (p_58_48 & g_47_32);
 assign p_58_48 = p_58_56 & p_55_48;
 assign g_58_48 = g_58_56 | (p_58_56 & g_55_48);
 assign p_58_56 = p_58_58 & p_57_56;
 assign g_58_56 = g_58_58 | (p_58_58 & g_57_56);
 assign sum[58] = p_58_58^ g_57_0;
 assign p_59_0 = p_59_32 & p_31_0;
 assign g_59_0 = g_59_32 | (p_59_32 & g_31_0);
 assign p_59_32 = p_59_48 & p_47_32;
 assign g_59_32 = g_59_48 | (p_59_48 & g_47_32);
 assign p_59_48 = p_59_56 & p_55_48;
 assign g_59_48 = g_59_56 | (p_59_56 & g_55_48);
 assign p_59_56 = p_59_58 & p_57_56;
 assign g_59_56 = g_59_58 | (p_59_58 & g_57_56);
 assign p_59_58 = p_59_59 & p_58_58;
 assign g_59_58 = g_59_59 | (p_59_59 & g_58_58);
 assign sum[59] = p_59_59^ g_58_0;
 assign p_60_0 = p_60_32 & p_31_0;
 assign g_60_0 = g_60_32 | (p_60_32 & g_31_0);
 assign p_60_32 = p_60_48 & p_47_32;
 assign g_60_32 = g_60_48 | (p_60_48 & g_47_32);
 assign p_60_48 = p_60_56 & p_55_48;
 assign g_60_48 = g_60_56 | (p_60_56 & g_55_48);
 assign p_60_56 = p_60_60 & p_59_56;
 assign g_60_56 = g_60_60 | (p_60_60 & g_59_56);
 assign sum[60] = p_60_60^ g_59_0;
 assign p_61_0 = p_61_32 & p_31_0;
 assign g_61_0 = g_61_32 | (p_61_32 & g_31_0);
 assign p_61_32 = p_61_48 & p_47_32;
 assign g_61_32 = g_61_48 | (p_61_48 & g_47_32);
 assign p_61_48 = p_61_56 & p_55_48;
 assign g_61_48 = g_61_56 | (p_61_56 & g_55_48);
 assign p_61_56 = p_61_60 & p_59_56;
 assign g_61_56 = g_61_60 | (p_61_60 & g_59_56);
 assign p_61_60 = p_61_61 & p_60_60;
 assign g_61_60 = g_61_61 | (p_61_61 & g_60_60);
 assign sum[61] = p_61_61^ g_60_0;
 assign p_62_0 = p_62_32 & p_31_0;
 assign g_62_0 = g_62_32 | (p_62_32 & g_31_0);
 assign p_62_32 = p_62_48 & p_47_32;
 assign g_62_32 = g_62_48 | (p_62_48 & g_47_32);
 assign p_62_48 = p_62_56 & p_55_48;
 assign g_62_48 = g_62_56 | (p_62_56 & g_55_48);
 assign p_62_56 = p_62_60 & p_59_56;
 assign g_62_56 = g_62_60 | (p_62_60 & g_59_56);
 assign p_62_60 = p_62_62 & p_61_60;
 assign g_62_60 = g_62_62 | (p_62_62 & g_61_60);
 assign sum[62] = p_62_62^ g_61_0;
 assign cout = g_62_0;
endmodule
